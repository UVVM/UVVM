-- This copy of OSVVM (UVVM OSVVM) has been modified in order to use the UVVM Utility Library.
--
-- Please see CHANGES.TXT for more information on the changes to the original OSVVM implementation.
-- Please see HOWTO-GUIDE.TXT for more information on how to use this copy of UVVM OSVVM.
--
--  Maintainer:        Bitvis AS     email:  support@bitvis.no
-- 

--
--  File Name:         OsvvmContext.vhd
--  Design Unit Name:  OsvvmContext
--  Revision:          STANDARD VERSION,  revision 2015.01
--
--  Maintainer:        Jim Lewis      email:  jim@synthworks.com--
--
--  Description
--      Context Declaration for OSVVM packages
--
--  Developed by/for:
--        SynthWorks Design Inc.
--        VHDL Training Classes
--        11898 SW 128th Ave.  Tigard, Or  97223
--        http://www.SynthWorks.com
--
--  Latest standard version available at:
--        http://www.SynthWorks.com/downloads
--
--  Revision History:      
--    Date      Version    Description
--    01/2015   2015.01    Initial Revision
--    06/2015   205.06     Added MemoryPkg
--
--
--  Copyright (c) 2015 by SynthWorks Design Inc.  All rights reserved.
--
--  Verbatim copies of this source file may be used and
--  distributed without restriction.
--
--  This source file is free software; you can redistribute it
--  and/or modify it under the terms of the ARTISTIC License
--  as published by The Perl Foundation; either version 2.0 of
--  the License, or (at your option) any later version.
--
--  This source is distributed in the hope that it will be
--  useful, but WITHOUT ANY WARRANTY; without even the implied
--  warranty of MERCHANTABILITY or FITNESS FOR A PARTICULAR
--  PURPOSE. See the Artistic License for details.
--
--  You should have received a copy of the license with this source.
--  If not download it from,
--     http://www.perlfoundation.org/artistic_license_2_0
--
--

context OsvvmContext is
    library uvvm_osvvm;  

    use uvvm_osvvm.NamePkg.all ;
    use uvvm_osvvm.TranscriptPkg.all ; 
    use uvvm_osvvm.OsvvmGlobalPkg.all ;
    use uvvm_osvvm.AlertLogPkg.all ; 
    use uvvm_osvvm.RandomPkg.all ;
    use uvvm_osvvm.CoveragePkg.all ;
    use uvvm_osvvm.MemoryPkg.all ;
    
end context OsvvmContext ; 

