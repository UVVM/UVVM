--========================================================================================================================
-- Copyright (c) 2018 by Bitvis AS.  All rights reserved.
-- You should have received a copy of the license file containing the MIT License (see LICENSE.TXT), if not,
-- contact Bitvis AS <support@bitvis.no>.
--
-- UVVM AND ANY PART THEREOF ARE PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND, EXPRESS OR IMPLIED, INCLUDING BUT NOT LIMITED TO THE
-- WARRANTIES OF MERCHANTABILITY, FITNESS FOR A PARTICULAR PURPOSE AND NONINFRINGEMENT. IN NO EVENT SHALL THE AUTHORS
-- OR COPYRIGHT HOLDERS BE LIABLE FOR ANY CLAIM, DAMAGES OR OTHER LIABILITY, WHETHER IN AN ACTION OF CONTRACT, TORT OR
-- OTHERWISE, ARISING FROM, OUT OF OR IN CONNECTION WITH UVVM OR THE USE OR OTHER DEALINGS IN UVVM.
--========================================================================================================================

------------------------------------------------------------------------------------------
-- Description   : See library quick reference (under 'doc') and README-file(s)
------------------------------------------------------------------------------------------

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

library uvvm_util;
context uvvm_util.uvvm_util_context;

use std.textio.all;

use work.csv_file_reader_pkg.all;
use work.local_adaptations_pkg.all;


package spec_cov_pkg is  


  alias config is shared_spec_cov_config;

  file RESULT_FILE : text;


  procedure initialize_req_cov(
    constant testcase         : string;
    constant req_list_file    : string;
    constant partial_cov_file : string
  );
  -- Overloading procedure, no req_list_file
  procedure initialize_req_cov(
    constant testcase         : string;
    constant partial_cov_file : string
  );


  procedure log_req_cov(
    constant requirement : string;
    constant testcase    : string;
    constant test_status : t_test_status  := NA;
    constant msg         : string         := "";
    constant scope       : string         := C_SCOPE
  );
  procedure log_req_cov(
    constant requirement : string;
    constant test_status : t_test_status  := NA;
    constant msg         : string         := "";
    constant scope       : string         := C_SCOPE
  );
  

  procedure finalize_req_cov(
    constant VOID : t_void
  );
  
  

  --=================================================================================================  
  -- Functions and procedures declared below this line are intended as internal functions
  --=================================================================================================  

  type t_line_vector is array(0 to config.max_testcases_per_req-1) of line;
  type t_requirement_entry is record
    valid         : boolean;
    requirement   : line;
    description   : line;
    num_tcs       : natural;
    tc_list       : t_line_vector;
  end record;
  type t_requirement_entry_array is array (natural range <>) of t_requirement_entry;

  -- Shared variables used internally in this context
  shared variable shared_csv_file               : csv_file_reader_type;
  shared variable shared_requirement_array      : t_requirement_entry_array(0 to config.max_testcases_per_req);
  shared variable shared_requirements_in_array  : natural := 0;

  constant C_FAIL_STRING                : string := "FAIL";
  constant C_PASS_STRING                : string := "PASS";

  procedure priv_log_entry(
    constant index : natural
  );

  procedure priv_read_and_parse_csv_file(
    constant req_list_file  : string
  );

  procedure priv_initialize_result_file(
    constant file_name : string
  );

  impure function priv_get_description(
    requirement : string;
    testcase    : string
  ) return string;

  impure function priv_requirement_exists(
    requirement : string
  ) return boolean;

  function priv_test_status_to_string(
    constant test_status : t_test_status
  ) return string;

  impure function priv_get_summary_string 
    return string;

  procedure priv_set_default_testcase_name(
    constant testcase : string
  );
  
  impure function priv_get_default_testcase_name 
  return string;

  impure function priv_find_string_length(
    constant search_string : string
  ) return natural;



end package spec_cov_pkg;


--=================================================================================================
--=================================================================================================
--=================================================================================================

package body spec_cov_pkg is

  -- private variables for pkg internal use only
  shared variable priv_testcase_name            : string(1 to C_CSV_FILE_MAX_LINE_LENGTH) := (others => NUL);
  shared variable priv_testcase_name_length     : natural;
  shared variable priv_testcase_passed          : boolean;
  shared variable priv_requirement_file_exists  : boolean;
  

  procedure initialize_req_cov(
    constant testcase         : string;
    constant req_list_file    : string;
    constant partial_cov_file : string
  ) is
  begin
    priv_set_default_testcase_name(testcase);
    -- update pkg local variables
    priv_testcase_passed          := true;
    priv_requirement_file_exists  := true;

    priv_read_and_parse_csv_file(req_list_file);    
    priv_initialize_result_file(partial_cov_file);
  end procedure initialize_req_cov;

  procedure initialize_req_cov(
    constant testcase         : string;
    constant partial_cov_file : string
  ) is
  begin
    log(ID_SPEC_COV, "Requirement Coverage initialized with no requirement file.", C_SCOPE);
    priv_set_default_testcase_name(testcase);
    -- update pkg local variables
    priv_testcase_passed          := true;
    priv_requirement_file_exists  := false;

    priv_initialize_result_file(partial_cov_file);
    end procedure initialize_req_cov;
  

  procedure log_req_cov(
    constant requirement : string;
    constant testcase    : string;
    constant test_status : t_test_status  := NA;
    constant msg         : string         := "";
    constant scope       : string         := C_SCOPE
  ) is
    variable v_requirement_to_file_line : line;
    variable v_requirement_status       : t_test_status := test_status;
  begin
    if shared_requirements_in_array = 0 and priv_requirement_file_exists = true then
      alert(TB_ERROR, "Requirements have not been parsed. Please used initialize_req_cov() with a requirement file before calling log_req_cov().", scope);
      return;
    end if;

    ---- Check if there were any errors globally
    if (shared_uvvm_status.found_unexpected_simulation_errors_or_worse = 1) then
      v_requirement_status := FAIL;
    end if;

    if v_requirement_status = FAIL then
      priv_testcase_passed := false;
    end if;

    -- Log result to transcript
    log(ID_SPEC_COV, "Logging requirement " & requirement & " [" & priv_test_status_to_string(v_requirement_status) & "]. '" & 
                      priv_get_description(requirement, testcase) & "'. " & msg, scope);

    -- Log to file
    write(v_requirement_to_file_line, requirement & C_CSV_DELIMITER & testcase & C_CSV_DELIMITER & priv_test_status_to_string(v_requirement_status));
    writeline(RESULT_FILE, v_requirement_to_file_line);
  end procedure log_req_cov;

  -- Overloading procedure
  procedure log_req_cov(
    constant requirement : string;
    constant test_status : t_test_status  := NA;
    constant msg         : string         := "";
    constant scope       : string         := C_SCOPE
  ) is 
  begin
    log_req_cov(requirement, priv_get_default_testcase_name , test_status, msg, scope);
  end procedure log_req_cov;
  
  
  procedure finalize_req_cov(
    constant VOID : t_void
  ) is
    variable v_checksum_string : line;
    constant c_summary_string  : string := priv_get_summary_string;
  begin
    -- Free used memory
    log(ID_SPEC_COV, "Freeing stored requirements from memory", C_SCOPE);

    for i in 0 to shared_requirements_in_array-1 loop
      deallocate(shared_requirement_array(i).requirement);
      deallocate(shared_requirement_array(i).description);
      for tc in 0 to shared_requirement_array(i).num_tcs-1 loop
        deallocate(shared_requirement_array(i).tc_list(tc));
      end loop;
      shared_requirement_array(i).num_tcs := 0;
      shared_requirement_array(i).valid   := false;
    end loop;
    shared_requirements_in_array := 0;
        
    -- Add closing line
    log(ID_SPEC_COV, "Marking requirement coverage result.", C_SCOPE);
    write(v_checksum_string, priv_get_summary_string);

    writeline(RESULT_FILE, v_checksum_string);

    file_close(RESULT_FILE);
    log(ID_SPEC_COV, "Requirement coverage finalized.", C_SCOPE);
  end procedure finalize_req_cov;
  


  
  --=================================================================================================  
  -- Functions and procedures declared below this line are intended as internal functions
  --=================================================================================================  


  procedure priv_initialize_result_file(
    constant file_name : string
  ) is
    variable v_file_open_status      : FILE_OPEN_STATUS;
    variable v_settings_to_file_line : line;
  
    constant c_note_string           : string := "NOTE: This coverage file is only valid when the last line is 'SUMMARY, " & 
                                                  priv_get_default_testcase_name & ", PASS'" & LF;
    constant c_testcase_string       : string := "TESTCASE_NAME: " & priv_get_default_testcase_name & LF;
    constant c_delimiter_string      : string := "DELIMITER: " & config.csv_delimiter & LF;
  begin
    file_open(v_file_open_status, RESULT_FILE, file_name, write_mode);
    check_file_open_status(v_file_open_status, file_name);

    -- Write setting to CSV file for Python script
    log(ID_SPEC_COV, "Adding test and configuration information to coverage file. ", C_SCOPE);
    write(v_settings_to_file_line, c_note_string);
    write(v_settings_to_file_line, c_testcase_string);
    write(v_settings_to_file_line, c_delimiter_string);
    writeline(RESULT_FILE, v_settings_to_file_line);
  end procedure priv_initialize_result_file;


  procedure priv_read_and_parse_csv_file(
      constant req_list_file  : string
  ) is 
    variable v_tc_valid : boolean;
    variable v_file_ok  : boolean;
  begin
    log(ID_SPEC_COV, "Reading and parsing requirement file, " & req_list_file, C_SCOPE);

    if shared_requirements_in_array > 0 then
      alert(TB_ERROR, "Requirements have already been read from file, please call finalize_req_cov before starting a new requirement coverage process.", C_SCOPE);
      return;
    end if;

    -- Open file and check status, return if failing
    v_file_ok := shared_csv_file.initialize(req_list_file, C_CSV_DELIMITER);
    if v_file_ok = false then
      return;
    end if;

    -- File ok, read file
    while not shared_csv_file.end_of_file loop
      shared_csv_file.readline;

      -- Read requirement
      shared_requirement_array(shared_requirements_in_array).requirement := new string'(shared_csv_file.read_string);
      -- Read description
      shared_requirement_array(shared_requirements_in_array).description := new string'(shared_csv_file.read_string);
      -- Read testcases
      v_tc_valid := true;
      shared_requirement_array(shared_requirements_in_array).num_tcs := 0;
      while v_tc_valid loop
        shared_requirement_array(shared_requirements_in_array).tc_list(shared_requirement_array(shared_requirements_in_array).num_tcs) := new string'(shared_csv_file.read_string);  
        if (shared_requirement_array(shared_requirements_in_array).tc_list(shared_requirement_array(shared_requirements_in_array).num_tcs).all(1) /= NUL) then
          shared_requirement_array(shared_requirements_in_array).num_tcs := shared_requirement_array(shared_requirements_in_array).num_tcs + 1;
        else
          v_tc_valid := false;
        end if;
      end loop;
      -- Validate entry
      shared_requirement_array(shared_requirements_in_array).valid := true;

      priv_log_entry(shared_requirements_in_array);
      shared_requirements_in_array := shared_requirements_in_array + 1;
    end loop;
        
    log(ID_SPEC_COV, "Closing requirement to testcase map file", C_SCOPE);
    shared_csv_file.dispose;
  end procedure priv_read_and_parse_csv_file;


  procedure priv_log_entry(
      constant index : natural
    ) is
  begin
    if shared_requirement_array(index).valid then
      -- log requirement and description to terminal
      log(ID_SPEC_COV, "Requirement: " & shared_requirement_array(index).requirement.all, C_SCOPE);
      log(ID_SPEC_COV, "Description: " & shared_requirement_array(index).description.all, C_SCOPE);
      -- log testcases to terminal
      for i in 0 to shared_requirement_array(index).num_tcs-1 loop
        log(ID_SPEC_COV, "  TC: " & shared_requirement_array(index).tc_list(i).all, C_SCOPE);
      end loop;
    else
      log(ID_SPEC_COV, "Requirement entry was not valid", C_SCOPE);
    end if;
  end procedure priv_log_entry;


  impure function priv_requirement_exists(
    requirement : string
  ) return boolean is
  begin
    for i in 0 to shared_requirements_in_array-1 loop
      if to_upper(shared_requirement_array(i).requirement.all(1 to requirement'length)) = to_upper(requirement(1 to requirement'length)) then
        return true;
      end if;
    end loop;
    return false;
  end function priv_requirement_exists;

  --impure function priv_requirement_and_tc_exists(
  --    requirement : string;
  --    testcase    : string
  --) return boolean is
  --begin
  --  for i in 0 to shared_requirements_in_array-1 loop
  --    if to_upper(shared_requirement_array(i).requirement.all(1 to requirement'length)) = to_upper(requirement(1 to requirement'length)) then
  --      for tc in 0 to shared_requirement_array(i).num_tcs-1 loop
  --        if to_upper(shared_requirement_array(i).tc_list(tc).all(1 to testcase'length)) = to_upper(testcase(1 to testcase'length)) then
  --          return true;
  --        end if;
  --      end loop;
  --    end if;
  --  end loop;
  --  return false;
  --end;

  impure function priv_get_description(
      requirement : string;
      testcase    : string
  ) return string is
  begin
    for i in 0 to shared_requirements_in_array-1 loop
      if shared_requirement_array(i).requirement.all(1 to requirement'length) = requirement(1 to requirement'length) then
        -- Found requirement
        for tc in 0 to shared_requirement_array(i).num_tcs-1 loop
          if shared_requirement_array(i).tc_list(tc).all(1 to testcase'length) = testcase(1 to testcase'length) then
            -- Found both requirement AND testcase
            return shared_requirement_array(i).description.all;
          end if;
        end loop;
      end if;
    end loop;

    if priv_requirement_file_exists = false then
      return "";
    else
      return "DESCRIPTION NOT FOUND";
    end if;
  end function priv_get_description;


  function priv_test_status_to_string(
    constant test_status : t_test_status
  ) return string is
  begin
    if test_status = PASS then
      return C_PASS_STRING;
    else -- test_status = FAIL
      return C_FAIL_STRING;
    end if;
  end function priv_test_status_to_string;


  impure function priv_get_summary_string 
    return string is
  begin
    -- Create a CSV coverage file summary string
    if (priv_testcase_passed = true) and (shared_uvvm_status.found_unexpected_simulation_errors_or_worse = 0) then
      return "SUMMARY, " & priv_get_default_testcase_name & ", " & C_PASS_STRING;
    else
      return "SUMMARY, " & priv_get_default_testcase_name & ", " & C_FAIL_STRING;
    end if;
  end function priv_get_summary_string;


  procedure priv_set_default_testcase_name(
    constant testcase : string
  ) is
  begin
    priv_testcase_name(1 to testcase'length)  := testcase;
  end procedure priv_set_default_testcase_name;


  impure function priv_get_default_testcase_name 
    return string is
    variable v_testcase_length : natural := priv_find_string_length(priv_testcase_name);
  begin 
    return priv_testcase_name(1 to v_testcase_length);
  end function priv_get_default_testcase_name;


  impure function priv_find_string_length(
    constant search_string : string
  ) return natural is
    variable v_return : natural := 0;
  begin
    -- loop string until NUL is found and return idx-1
    for idx in 1 to search_string'length loop
      if search_string(idx) = NUL then
        return idx - 1;
      end if;
    end loop;

    -- NUL was not found, return full length
    return search_string'length;
  end function priv_find_string_length;

end package body spec_cov_pkg;
