--================================================================================================================================
-- Copyright (c) 2020 by Bitvis AS.  All rights reserved.
-- You should have received a copy of the license file containing the MIT License (see LICENSE.TXT), if not,
-- contact Bitvis AS <support@bitvis.no>.
--
-- UVVM AND ANY PART THEREOF ARE PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND, EXPRESS OR IMPLIED, INCLUDING BUT NOT LIMITED TO
-- THE WARRANTIES OF MERCHANTABILITY, FITNESS FOR A PARTICULAR PURPOSE AND NONINFRINGEMENT. IN NO EVENT SHALL THE AUTHORS
-- OR COPYRIGHT HOLDERS BE LIABLE FOR ANY CLAIM, DAMAGES OR OTHER LIABILITY, WHETHER IN AN ACTION OF CONTRACT, TORT OR
-- OTHERWISE, ARISING FROM, OUT OF OR IN CONNECTION WITH UVVM OR THE USE OR OTHER DEALINGS IN UVVM.
--================================================================================================================================

---------------------------------------------------------------------------------------------
-- Description : See library quick reference (under 'doc') and README-file(s)
---------------------------------------------------------------------------------------------

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

library uvvm_util;
context uvvm_util.uvvm_util_context;

library uvvm_vvc_framework;
use uvvm_vvc_framework.ti_vvc_framework_support_pkg.all;

entity hvvc_to_vvc_bridge is
  generic(
    GC_INSTANCE_IDX        : integer;
    GC_DUT_IF_FIELD_CONFIG : t_dut_if_field_config_direction_array;
    GC_MAX_NUM_BYTES       : positive;
    GC_PHY_MAX_ACCESS_TIME : time;
    GC_SCOPE               : string
  );
  port(
    hvvc_to_bridge : in  t_hvvc_to_bridge(data_bytes(0 to GC_MAX_NUM_BYTES-1));
    bridge_to_hvvc : out t_bridge_to_hvvc(data_bytes(0 to GC_MAX_NUM_BYTES-1))
  );
end entity hvvc_to_vvc_bridge;