--================================================================================================================================
-- Copyright 2024 UVVM
-- Licensed under the Apache License, Version 2.0 (the "License"); you may not use this file except in compliance with the License.
-- You may obtain a copy of the License at http://www.apache.org/licenses/LICENSE-2.0 and in the provided LICENSE.TXT.
--
-- Unless required by applicable law or agreed to in writing, software distributed under the License is distributed on
-- an "AS IS" BASIS, WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
-- See the License for the specific language governing permissions and limitations under the License.
--================================================================================================================================
-- Note : Any functionality not explicitly described in the documentation is subject to change at any time
----------------------------------------------------------------------------------------------------------------------------------

------------------------------------------------------------------------------------------
-- Description   : See library quick reference (under 'doc') and README-file(s)
------------------------------------------------------------------------------------------

context vvc_framework_context is
  library uvvm_vvc_framework;
  use uvvm_vvc_framework.ti_data_fifo_pkg.all;
  use uvvm_vvc_framework.ti_data_queue_pkg.all;
  use uvvm_vvc_framework.ti_data_stack_pkg.all;
  use uvvm_vvc_framework.ti_vvc_framework_support_pkg.all;
  use uvvm_vvc_framework.ti_protected_types_pkg.all;
end context;