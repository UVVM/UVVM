-------------------------------------------------------
--  Copyright (c) 2011 Xilinx Inc.
--  All Right Reserved.
-------------------------------------------------------
--
--   ____  ____
--  /   /\/   / 
-- /___/  \  /     Vendor      : Xilinx 
-- \   \   \/      Version : 11.1
--  \   \          Description : 
--  /   /                      
-- /___/   /\      Filename    : BUFG_LB.vhd
-- \   \  /  \      
--  \__ \/\__ \                   
--                                 
--  Generated by    : /home/chen/xfoundry/HEAD/env/Databases/CAEInterfaces/LibraryWriters/bin/ltw.pl
--  Revision: 1.0
--    11/15/11 - 634082 - connected ouput.
--  End Revision
-------------------------------------------------------

----- CELL BUFG_LB -----

library IEEE;
use IEEE.STD_LOGIC_arith.all;
use IEEE.STD_LOGIC_1164.all;

library unisim;
use unisim.VCOMPONENTS.all;
use unisim.vpkg.all;

  entity BUFG_LB is
    port (
      CLKOUT               : out std_ulogic;
      CLKIN                : in std_ulogic      
    );
  end BUFG_LB;

  architecture BUFG_LB_V of BUFG_LB is
  begin
    
    CLKOUT <= TO_X01(CLKIN);

  end BUFG_LB_V;
