--========================================================================================================================
-- Copyright (c) 2016 by Bitvis AS.  All rights reserved.
-- You should have received a copy of the license file containing the MIT License (see LICENSE.TXT), if not, 
-- contact Bitvis AS <support@bitvis.no>.
--
-- UVVM AND ANY PART THEREOF ARE PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND, EXPRESS OR IMPLIED, INCLUDING BUT NOT LIMITED TO THE
-- WARRANTIES OF MERCHANTABILITY, FITNESS FOR A PARTICULAR PURPOSE AND NONINFRINGEMENT. IN NO EVENT SHALL THE AUTHORS
-- OR COPYRIGHT HOLDERS BE LIABLE FOR ANY CLAIM, DAMAGES OR OTHER LIABILITY, WHETHER IN AN ACTION OF CONTRACT, TORT OR
-- OTHERWISE, ARISING FROM, OUT OF OR IN CONNECTION WITH UVVM OR THE USE OR OTHER DEALINGS IN UVVM.
--========================================================================================================================

------------------------------------------------------------------------------------------
-- VHDL unit     : Bitvis AVALON_MM Library : avalon_mm_spi_tb
--
-- Description   : See dedicated powerpoint presentation and README-file(s)
------------------------------------------------------------------------------------------

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

library STD;
use std.textio.all;

library vunit_lib;
context vunit_lib.vunit_run_context;

library uvvm_util;
use uvvm_util.types_pkg.all;
use uvvm_util.string_methods_pkg.all;
use uvvm_util.adaptations_pkg.all;
use uvvm_util.methods_pkg.all;
use uvvm_util.bfm_common_pkg.all;

library bitvis_vip_avalon_mm;
use bitvis_vip_avalon_mm.avalon_mm_bfm_pkg.all;

-- Test case entity
entity avalon_mm_spi_tb is
  generic (
    -- This generic is used to configure the testbench from run.py, e.g. what
    -- test case to run. The default value is used when not running from script
    -- and in that case all test cases are run.
    runner_cfg : runner_cfg_t := runner_cfg_default);
end entity;

-- Test case architecture
architecture func of avalon_mm_spi_tb is

  constant C_CLK_PERIOD  : time := 10 ns;
  signal clk : std_logic;

  -- signals
  -- The avalon_mm interface is gathered in two records (to and from DUT), 
  -- so procedures that use the avalon_mm interface have less arguments
  signal avalon_mm_if : t_avalon_mm_if(address(2 downto 0), byte_enable(1 downto 0), writedata(15 downto 0), readdata(15 downto 0));
  signal clock_ena       : boolean := false;

  -- SPI signals
  signal MISO          :  STD_LOGIC;
  signal MOSI          :  STD_LOGIC;
  signal SCLK          :  STD_LOGIC;
  signal SS_n          :  STD_LOGIC;
  signal dataavailable :  STD_LOGIC;
  signal endofpacket   :  STD_LOGIC;
  signal irq           :  STD_LOGIC;
  signal readyfordata  :  STD_LOGIC;
  
  component avalon_spi
    port (
      signal MISO          : IN  STD_LOGIC;
      signal clk           : IN  STD_LOGIC;
      signal data_from_cpu : IN  STD_LOGIC_VECTOR (15 DOWNTO 0);
      signal mem_addr      : IN  STD_LOGIC_VECTOR (2 DOWNTO 0);
      signal read_n        : IN  STD_LOGIC;
      signal reset_n       : IN  STD_LOGIC;
      signal spi_select    : IN  STD_LOGIC;
      signal write_n       : IN  STD_LOGIC;
      signal MOSI          : OUT STD_LOGIC;
      signal SCLK          : OUT STD_LOGIC;
      signal SS_n          : OUT STD_LOGIC;
      signal data_to_cpu   : OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
      signal dataavailable : OUT STD_LOGIC;
      signal endofpacket   : OUT STD_LOGIC;
      signal irq           : OUT STD_LOGIC;
      signal readyfordata  : OUT STD_LOGIC);
  end component;
begin

  -- Set up clock generator
  p_clock: clock_generator(clk, clock_ena, C_CLK_PERIOD, "Avalon MM clock");

  -----------------------------------------------------------------------------
  -- Instantiate DUT - a master mode Avalon_Mm SPI
  -----------------------------------------------------------------------------
  avalon_spi_1: avalon_spi
    port map (
      MISO          => MISO,
      clk           => clk,
      data_from_cpu => avalon_mm_if.writedata(15 downto 0),
      mem_addr      => avalon_mm_if.address(2 downto 0),
      read_n        => not avalon_mm_if.read,
      reset_n       => not avalon_mm_if.reset,
      spi_select    => avalon_mm_if.chipselect,
      write_n       => not avalon_mm_if.write,
      MOSI          => MOSI,
      SCLK          => SCLK,
      SS_n          => SS_n,
      data_to_cpu   => avalon_mm_if.readdata(15 downto 0),
      dataavailable => dataavailable,
      endofpacket   => endofpacket,
      irq           => irq,
      readyfordata  => readyfordata);
      
  -- Response signal is not used in the DUT, so we ground it.
  avalon_mm_if.response <= (others => '0');

  p_loopback_mosi: process (MOSI)
  begin  -- process MOSI
    MISO <= MOSI;
  end process p_loopback_mosi;
  ------------------------------------------------
  -- PROCESS: p_main
  ------------------------------------------------
  p_main: process
    constant C_SCOPE     : string  := C_TB_SCOPE_DEFAULT;
    -- BFM config
    variable avalon_mm_bfm_config : t_avalon_mm_bfm_config := C_avalon_mm_bfm_config_DEFAULT;

    -- Overloads for simplification
    procedure log(
      msg   : string) is
    begin
      log(ID_SEQUENCER, msg, C_SCOPE);
    end;

    -- overload for this testbench
    procedure avalon_mm_write (
      addr_value           : in unsigned;
      data_value           : in std_logic_vector;
      alert_level          : in t_alert_level := error
      ) is
      variable timeout : boolean := false;
      variable cycle   : natural := 0;
    begin
      if addr_value = 1 then
        -- check that SPI module is ready for data - wait if necessary
        while not readyfordata loop
          wait until rising_edge(clk);
          cycle := cycle+1;
          if cycle = 100 then
            timeout := true;
            alert(alert_level, "avalon_mm_write() timeout waiting for SPI to be ready");
            exit;
          end if;
        end loop;
        if not timeout then
          avalon_mm_write(addr_value, data_value, "", clk, avalon_mm_if, "11", C_SCOPE, shared_msg_id_panel, avalon_mm_bfm_config);
        end if;
      else
        avalon_mm_write(addr_value, data_value, "", clk, avalon_mm_if, "11", C_SCOPE, shared_msg_id_panel, avalon_mm_bfm_config);
      end if;
    end;
    
    -- overload for this testbench
    procedure avalon_mm_read (
      addr_value           : in unsigned;
      data_value           : out std_logic_vector;
      alert_level          : in t_alert_level := error
      ) is
      variable timeout : boolean := false;
      variable cycle   : natural := 0;
    begin
      if addr_value = 0 then
        -- check that SPI module is ready to deliver - wait if necessary
        while not dataavailable loop
          wait until rising_edge(clk);
          cycle := cycle+1;
          if cycle = 100 then
            timeout := true;
            alert(alert_level, "avalon_mm_read) timeout waiting for SPI to have data");
            exit;
          end if;
        end loop;
        if not timeout then
          avalon_mm_read(addr_value, data_value, "", clk, avalon_mm_if, C_SCOPE, shared_msg_id_panel, avalon_mm_bfm_config);
        end if;
      else
        avalon_mm_read(addr_value, data_value, "", clk, avalon_mm_if, C_SCOPE, shared_msg_id_panel, avalon_mm_bfm_config);
      end if;
    end;

    -- overload for this testbench
    procedure avalon_mm_check (
      addr_value           : in unsigned;
      data_exp             : in std_logic_vector;
      alert_level          : in t_alert_level := error
      ) is
      variable timeout : boolean := false;
      variable cycle   : natural := 0;
    begin
      -- same timeout as for reads - if checking addr 0
      if addr_value = 0 then
        -- check that SPI module is ready to deliver - wait if necessary
        while not dataavailable loop
          wait until rising_edge(clk);
          cycle := cycle+1;
          if cycle = 100 then
            timeout := true;
            alert(alert_level, "avalon_mm_read) timeout waiting for SPI to have data");
            exit;
          end if;
        end loop;
        if not timeout then
          avalon_mm_check(addr_value, data_exp, "", clk, avalon_mm_if, alert_level, C_SCOPE, shared_msg_id_panel, avalon_mm_bfm_config);
        end if;
      else
        avalon_mm_check(addr_value, data_exp, "", clk, avalon_mm_if, alert_level, C_SCOPE, shared_msg_id_panel, avalon_mm_bfm_config);
      end if;
    end;
    
    variable i              : integer;
    variable fifo_data       : std_logic_vector(31 downto 0);
    variable v_alert_num_mismatch : boolean := false;

  begin
    
    -- To avoid that log files from different test cases (run in separate
    -- simulations) overwrite each other run.py provides separate test case
    -- directories through the runner_cfg generic (<root>/vunit_out/tests/<test case
    -- name>). When not using run.py the default path is the current directory
    -- (<root>/vunit_out/<simulator>). These directories are used by VUnit
    -- itself and these lines make sure that BVUL do to.
    set_log_file_name(join(output_path(runner_cfg), "_Log.txt"));
    set_alert_file_name(join(output_path(runner_cfg), "_Alert.txt"));
    
    -- Setup the VUnit runner with the input configuration.
    test_runner_setup(runner, runner_cfg);
    
    -- The default behavior for VUnit is to stop the simulation on a failing
    -- check when running from script but keep on running when running without
    -- script. The rationale for this and how you can change that behavior is
    -- described at the bottom of this file (see Stopping the Simulation on
    -- Failing Checks). The following if statement causes BVUL checks to behave
    -- in the same way.
    if not active_python_runner(runner_cfg) then
      set_alert_stop_limit(ERROR, 0);
    end if;
  
    -- set up our avalon_mm config - could be different than default config in BFM
    avalon_mm_bfm_config.clock_period             := C_CLK_PERIOD;  -- same clock period for BFM as for clock generator
    avalon_mm_bfm_config.max_wait_cycles          := 10;
    avalon_mm_bfm_config.num_wait_states          := 1;
    avalon_mm_bfm_config.use_waitrequest          := false;
    avalon_mm_bfm_config.use_readdatavalid        := false;
    
    -- Print the configuration to the log
    report_global_ctrl(VOID);
    report_msg_id_panel(VOID);

    enable_log_msg(ALL_MESSAGES);
    --disable_log_msg(ALL_MESSAGES);
    --enable_log_msg(ID_LOG_HDR);

    log("Start Simulation of TB for AVALON_MM");
    ------------------------------------------------------------
    clock_ena <= true; -- the avalon_mm_reset routine assumes the clock is running
    avalon_mm_reset(clk, avalon_mm_if, 5, "Resetting Avalon MM Interface", C_SCOPE, shared_msg_id_panel, avalon_mm_bfm_config);

    -- allow some time before we start
    for i in 0 to 50 loop
      wait until rising_edge(clk);
    end loop;
    
    log("Write to TXDATA register");
    avalon_mm_write("1", x"55");
    avalon_mm_write("1", x"aa");

    -- should take 8 bits X 10 clocks (SPI clock 10 x slower)
    for i in 0 to 80 loop
      wait until rising_edge(clk);
    end loop;
    
    log("Read back (and check) loopback of TXDATA");
    avalon_mm_check("0", x"55");
    avalon_mm_check("0", x"aa");
    
    --==================================================================================================
    -- Ending the simulation
    --------------------------------------------------------------------------------------
    -- allow some time for completion
    for i in 0 to 100 loop
      wait until rising_edge(clk);
    end loop;
    
    report_alert_counters(VOID); -- Report final counters and print conclusion for simulation (Success/Fail)
    log("SIMULATION COMPLETED");
    
    -- Cleanup VUnit. The UVVM-Util error status is imported into VUnit at this
    -- point. This is neccessary when the UVVM-Util alert stop limit is set such that
    -- UVVM-Util doesn't stop on the first error. In that case VUnit has no way of
    -- knowing the error status unless you tell it.
    for alert_level in NOTE to t_alert_level'right loop
      if alert_level /= MANUAL_CHECK and get_alert_counter(alert_level, REGARD) /= get_alert_counter(alert_level, EXPECT) then
        v_alert_num_mismatch := true;
      end if;
    end loop;
    
    test_runner_cleanup(runner, v_alert_num_mismatch);
    wait;

  end process p_main;

end func;
