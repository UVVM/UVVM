--========================================================================================================================
-- Copyright (c) 2017 by Bitvis AS.  All rights reserved.
-- You should have received a copy of the license file containing the MIT License (see LICENSE.TXT), if not,
-- contact Bitvis AS <support@bitvis.no>.
--
-- UVVM AND ANY PART THEREOF ARE PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND, EXPRESS OR IMPLIED, INCLUDING BUT NOT LIMITED TO THE
-- WARRANTIES OF MERCHANTABILITY, FITNESS FOR A PARTICULAR PURPOSE AND NONINFRINGEMENT. IN NO EVENT SHALL THE AUTHORS
-- OR COPYRIGHT HOLDERS BE LIABLE FOR ANY CLAIM, DAMAGES OR OTHER LIABILITY, WHETHER IN AN ACTION OF CONTRACT, TORT OR
-- OTHERWISE, ARISING FROM, OUT OF OR IN CONNECTION WITH UVVM OR THE USE OR OTHER DEALINGS IN UVVM.
--========================================================================================================================

------------------------------------------------------------------------------------------
-- Description   : See library quick reference (under 'doc') and README-file(s)
------------------------------------------------------------------------------------------

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

library vunit_lib;
context vunit_lib.vunit_run_context;

library uvvm_util;
context uvvm_util.uvvm_util_context;

library uvvm_vvc_framework;
use uvvm_vvc_framework.ti_vvc_framework_support_pkg.all;

library bitvis_vip_sbi;
context bitvis_vip_sbi.vvc_context;
use bitvis_vip_sbi.sbi_bfm_pkg.all;


-- Test case entity
entity sbi_tb is
  generic (
    -- This generic is used to configure the testbench from run.py, e.g. what
    -- test case to run. The default value is used when not running from script
    -- and in that case all test cases are run.
    runner_cfg : runner_cfg_t := runner_cfg_default);
end entity;

-- Test case architecture
architecture func of sbi_tb is

  constant C_CLK_PERIOD   : time := 10 ns;    -- **** Trenger metode for setting av clk period
  constant C_SCOPE        : string := "SBI_VVC_TB";

  -- FIFO Register map :
  constant C_ADDR_FIFO_PUT            : unsigned := "000";
  constant C_ADDR_FIFO_GET            : unsigned := "001";
  constant C_ADDR_FIFO_COUNT          : unsigned := "010";
  constant C_ADDR_FIFO_PEEK           : unsigned := "011";
  constant C_ADDR_FIFO_FLUSH          : unsigned := "100";
  constant C_ADDR_FIFO_MAX_COUNT      : unsigned := "101";
  constant C_DATA_DONTCARE            : std_logic_vector(7 downto 0) := x"00";


begin

  -----------------------------------------------------------------------------
  -- Instantiate test harness, containing DUT and Executors
  -----------------------------------------------------------------------------
  i_test_harness : entity work.test_harness generic map(GC_CLK_PERIOD => C_CLK_PERIOD);

  i_ti_uvvm_engine  : entity uvvm_vvc_framework.ti_uvvm_engine;


  ------------------------------------------------
  -- PROCESS: p_main
  ------------------------------------------------
  p_main: process

      -- BFM config
      variable sbi_bfm_config       : t_sbi_bfm_config := C_SBI_BFM_CONFIG_DEFAULT;

      variable v_cmd_idx            : integer;
      variable v_data               : work.vvc_cmd_pkg.t_vvc_result;
      variable v_is_ok              : boolean := false;
      variable v_timestamp          : time;
      variable v_alert_num_mismatch : boolean := false;

      alias clk     is << signal i_test_harness.clk      : std_logic >>;
      alias sbi1_if is << signal i_test_harness.sbi_if_1 : t_sbi_if >>;

  begin

    -- To avoid that log files from different test cases (run in separate
    -- simulations) overwrite each other run.py provides separate test case
    -- directories through the runner_cfg generic (<root>/vunit_out/tests/<test case
    -- name>). When not using run.py the default path is the current directory
    -- (<root>/vunit_out/<simulator>). These directories are used by VUnit
    -- itself and these lines make sure that BVUL do to.
    set_log_file_name(join(output_path(runner_cfg), "_Log.txt"));
    set_alert_file_name(join(output_path(runner_cfg), "_Alert.txt"));

    -- Setup the VUnit runner with the input configuration.
    test_runner_setup(runner, runner_cfg);



    -- The default behavior for VUnit is to stop the simulation on a failing
    -- check when running from script but keep on running when running without
    -- script. The rationale for this and how you can change that behavior is
    -- described at the bottom of this file (see Stopping the Simulation on
    -- Failing Checks). The following if statement causes BVUL checks to behave
    -- in the same way.
    if not active_python_runner(runner_cfg) then
      set_alert_stop_limit(ERROR, 0);
    end if;

    await_uvvm_initialization(VOID);

    set_alert_stop_limit(TB_ERROR,4);

    disable_log_msg(ALL_MESSAGES);
    enable_log_msg(ID_SEQUENCER);
    enable_log_msg(ID_LOG_HDR);
    enable_log_msg(ID_BFM);
    enable_log_msg(ID_BFM_POLL);

    disable_log_msg(VVC_BROADCAST, ALL_MESSAGES);
    enable_log_msg(VVC_BROADCAST, ID_BFM);
    enable_log_msg(VVC_BROADCAST, ID_BFM_POLL);

    --disable_log_msg(SBI_VVCT, 1, ALL_MESSAGES);
    --enable_log_msg(SBI_VVCT, 1, ID_BFM);
    --enable_log_msg(SBI_VVCT, 1, ID_BFM_POLL);
    --
    --disable_log_msg(SBI_VVCT, 2, ALL_MESSAGES);
    --enable_log_msg(SBI_VVCT, 2, ID_BFM);
    --enable_log_msg(SBI_VVCT, 2, ID_BFM_POLL);

    -- Print the configuration to the log
    report_global_ctrl(VOID);
    report_msg_id_panel(VOID);

    -- Set that ready signal is not in use
    shared_sbi_vvc_config(1).bfm_config.use_ready_signal := false;
    shared_sbi_vvc_config(2).bfm_config.use_ready_signal := false;

    sbi_bfm_config.clock_period         := C_CLK_PERIOD;
    sbi_bfm_config.setup_time           := C_CLK_PERIOD/4;
    sbi_bfm_config.hold_time            := C_CLK_PERIOD/4;
    wait for 3*C_CLK_PERIOD;  -- Wait for reset being released in test harness

    while test_suite loop
      --------------------------------------------------------------------------------------
      -- Verifying
      --------------------------------------------------------------------------------------
      if run("simple_write_and_check") then
        log(ID_LOG_HDR, "Test of simple write and check", C_SCOPE);
        --==========================================================================

        log("Write with both interfaces");
        sbi_write(SBI_VVCT,1, C_ADDR_FIFO_PUT, x"AA", "Write PUT on FIFO 1");
        sbi_write(SBI_VVCT,2, C_ADDR_FIFO_PUT, x"FF", "Write PUT on FIFO 2");
        await_completion(SBI_VVCT,1, 16 ns, "Await execution");

        log("Read and check with both interfaces");
        sbi_check(SBI_VVCT,1, C_ADDR_FIFO_GET, x"FF", "Check GET data on FIFO 2", ERROR);
        sbi_check(SBI_VVCT,2, C_ADDR_FIFO_GET, x"AA", "Check GET data on FIFO 1", ERROR);
        await_completion(SBI_VVCT,1, 16 ns, "Await execution");

    elsif run("simple_write_and_read") then
        log(ID_LOG_HDR, "Test of simple write and read", C_SCOPE);
        --==========================================================================
        -- Write to FIFO
        log("Write with both interfaces");
        sbi_write(SBI_VVCT,1, C_ADDR_FIFO_PUT, x"12", "Write PUT on FIFO 1");
        sbi_write(SBI_VVCT,2, C_ADDR_FIFO_PUT, x"53", "Write PUT on FIFO 2");
        await_completion(SBI_VVCT,1, 16 ns, "Await execution");

        -- Read, fetch and check on FIFO 2
        log("Read and check FIFO 2 using SBI IF 1");
        sbi_read(SBI_VVCT,1, C_ADDR_FIFO_GET, "Read from FIFO 2 and store result in VVC");
        v_cmd_idx := get_last_received_cmd_idx(SBI_VVCT, 1); -- for last read
        await_completion(SBI_VVCT,1, v_cmd_idx, 100 ns, "Wait for sbi_read to finish");
        fetch_result(SBI_VVCT,1, v_cmd_idx, v_data, v_is_ok,  "Fetching read-result");
        check_value(v_is_ok, ERROR, "Readback OK via fetch_result()");
        check_value(v_data(7 downto 0), x"53", ERROR, "Readback data via fetch_result()");

        -- Read, fetch and check on FIFO 1
        log("Read and check FIFO 1 using SBI IF 2");
        sbi_read(SBI_VVCT,2, C_ADDR_FIFO_GET, "Read from FIFO 1 and store result in VVC");
        v_cmd_idx := get_last_received_cmd_idx(SBI_VVCT, 2); -- for last read
        await_completion(SBI_VVCT,2, v_cmd_idx, 100 ns, "Wait for sbi_read to finish");
        fetch_result(SBI_VVCT,2, v_cmd_idx, v_data, v_is_ok, "Fetching read-result");
        check_value(v_is_ok, ERROR, "Readback OK via fetch_result()");
        check_value(v_data(7 downto 0), x"12", ERROR, "Readback data via fetch_result()");

        await_completion(SBI_VVCT,2, 100 ns, "Await execution");

    elsif run("test_of_poll_until") then
        log(ID_LOG_HDR, "Test of poll until", C_SCOPE);
        --==========================================================================

        -- Fill FIFO 1
        sbi_write(SBI_VVCT,1, C_ADDR_FIFO_PUT, x"01", "Write PUT on FIFO 1");
        sbi_write(SBI_VVCT,1, C_ADDR_FIFO_PUT, x"56", "Write PUT on FIFO 1");
        sbi_write(SBI_VVCT,1, C_ADDR_FIFO_PUT, x"a3", "Write PUT on FIFO 1");
        sbi_write(SBI_VVCT,1, C_ADDR_FIFO_PUT, x"4d", "Write PUT on FIFO 1");
        sbi_write(SBI_VVCT,1, C_ADDR_FIFO_PUT, x"00", "Write PUT on FIFO 1");
        sbi_write(SBI_VVCT,1, C_ADDR_FIFO_PUT, x"42", "Write PUT on FIFO 1");
        await_completion(SBI_VVCT,1, 1000 ns, "Await execution");

        -- Fill FIFO 2
        sbi_write(SBI_VVCT,2, C_ADDR_FIFO_PUT, x"01", "Write PUT on FIFO 2");
        sbi_write(SBI_VVCT,2, C_ADDR_FIFO_PUT, x"56", "Write PUT on FIFO 2");
        sbi_write(SBI_VVCT,2, C_ADDR_FIFO_PUT, x"a3", "Write PUT on FIFO 2");
        sbi_write(SBI_VVCT,2, C_ADDR_FIFO_PUT, x"4d", "Write PUT on FIFO 2");
        sbi_write(SBI_VVCT,2, C_ADDR_FIFO_PUT, x"00", "Write PUT on FIFO 2");
        sbi_write(SBI_VVCT,2, C_ADDR_FIFO_PUT, x"42", "Write PUT on FIFO 2");
        await_completion(SBI_VVCT,2, 1000 ns, "Await execution");

        -- Poll from FIFO 2
        sbi_poll_until(SBI_VVCT,1, C_ADDR_FIFO_GET,  x"42", "Test of POLL_UNTIL within 100 ns", 0, 100 ns, ERROR);

        -- Poll from FIFO 1
        sbi_poll_until(SBI_VVCT,2, C_ADDR_FIFO_GET,  x"42", "Test of POLL_UNTIL within 10 occurrences", 10, 0 ns, ERROR);

        await_completion(SBI_VVCT,1, 1000 ns, "Await execution");
        await_completion(SBI_VVCT,2, 1000 ns, "Await execution");

      elsif run("extended_write_and_read") then
        log(ID_LOG_HDR, "Test of write and read from other addresses on both VVCs", C_SCOPE);
        --==========================================================================

        sbi_write(SBI_VVCT,1, C_ADDR_FIFO_FLUSH, C_DATA_DONTCARE, "Flush FIFO 1");
        sbi_write(SBI_VVCT,2, C_ADDR_FIFO_FLUSH, C_DATA_DONTCARE, "Flush FIFO 2");

        sbi_check(SBI_VVCT,2, C_ADDR_FIFO_COUNT, x"00", "Check that FIFO 1 is empty", ERROR);
        sbi_check(SBI_VVCT,1, C_ADDR_FIFO_COUNT, x"00", "Check that FIFO 2 is empty", ERROR);

        sbi_write(SBI_VVCT,1, C_ADDR_FIFO_PUT, x"11", "Write PUT on FIFO 1");
        sbi_write(SBI_VVCT,1, C_ADDR_FIFO_PUT, x"12", "Write PUT on FIFO 1");
        sbi_write(SBI_VVCT,1, C_ADDR_FIFO_PUT, x"13", "Write PUT on FIFO 1");
        sbi_write(SBI_VVCT,2, C_ADDR_FIFO_PUT, x"11", "Write PUT on FIFO 2");
        sbi_write(SBI_VVCT,2, C_ADDR_FIFO_PUT, x"12", "Write PUT on FIFO 2");
        sbi_write(SBI_VVCT,2, C_ADDR_FIFO_PUT, x"13", "Write PUT on FIFO 2");

        sbi_check(SBI_VVCT,2, C_ADDR_FIFO_COUNT, x"18", "Check that FIFO 1 has three elements (3*8bit = 24 = x'18')", ERROR);
        sbi_check(SBI_VVCT,1, C_ADDR_FIFO_COUNT, x"18", "Check that FIFO 2 has three elements (3*8bit = 24 = x'18')", ERROR);

        sbi_check(SBI_VVCT,2, C_ADDR_FIFO_PEEK, x"11", "Peek on FIFO 1", ERROR);
        sbi_check(SBI_VVCT,2, C_ADDR_FIFO_PEEK, x"11", "Peek on FIFO 1 again", ERROR);
        sbi_check(SBI_VVCT,1, C_ADDR_FIFO_PEEK, x"11", "Peek on FIFO 2", ERROR);
        sbi_check(SBI_VVCT,1, C_ADDR_FIFO_PEEK, x"11", "Peek on FIFO 2 again", ERROR);

        sbi_write(SBI_VVCT,1, C_ADDR_FIFO_FLUSH, C_DATA_DONTCARE, "Flush FIFO 1");
        sbi_write(SBI_VVCT,2, C_ADDR_FIFO_FLUSH, C_DATA_DONTCARE, "Flush FIFO 2");

        sbi_check(SBI_VVCT,2, C_ADDR_FIFO_COUNT, x"00", "Check that FIFO 1 is empty", ERROR);
        sbi_check(SBI_VVCT,1, C_ADDR_FIFO_COUNT, x"00", "Check that FIFO 2 is empty", ERROR);

        await_completion(SBI_VVCT,1, 1000 ns, "Await execution");
        await_completion(SBI_VVCT,2, 1000 ns, "Await execution");

      elsif run("read_of_previous_value") then
        -- Test DIVERSE
        log(ID_LOG_HDR, "Test read of a previous value");
        ------------------------------------------------------
        sbi_write(SBI_VVCT,1, C_ADDR_FIFO_PUT, x"A0", "Write PUT on FIFO 1");
        sbi_write(SBI_VVCT,1, C_ADDR_FIFO_PUT, x"B1", "Write PUT on FIFO 1");
        sbi_write(SBI_VVCT,1, C_ADDR_FIFO_PUT, x"C2", "Write PUT on FIFO 1");
        await_completion(SBI_VVCT, 1, 100 ns);

        log("\rNow starting readback with 100T delay between 1st and 2nd read");
        sbi_read(SBI_VVCT,2, C_ADDR_FIFO_GET, "Readback inside VVC");
        v_cmd_idx := get_last_received_cmd_idx(SBI_VVCT, 2); -- for last read
        insert_delay(SBI_VVCT,2, 100, "100T delay");
        sbi_read(SBI_VVCT,2, C_ADDR_FIFO_GET, "Readback inside VVC");
        sbi_read(SBI_VVCT,2, C_ADDR_FIFO_GET, "Readback inside VVC");
        v_timestamp := now;

        log("\rFetch the 1st result");
        await_completion(SBI_VVCT,2, v_cmd_idx, 100 ns, "first read should be executed immediately");
        fetch_result(SBI_VVCT,2, v_cmd_idx, v_data, v_is_ok, "Fetching available read-result");
        check_value(v_is_ok, ERROR, "Readback OK via fetch_result()");
        check_value(v_data(7 downto 0), x"A0", ERROR, "Readback data via fetch_result()");

        log("\rFetch the 2nd result");
        await_completion(SBI_VVCT,2, v_cmd_idx+2, 110 * C_CLK_PERIOD, "2nd read should be executed 100 cycles after the first");
        fetch_result(SBI_VVCT,2, v_cmd_idx+2, v_data, v_is_ok, "Fetching 2nd read-result");
        check_value(v_is_ok, ERROR, "Readback OK via fetch_result()");
        check_value(v_data(7 downto 0), x"B1", ERROR, "Readback data via fetch_result()");
        check_value_in_range((now-v_timestamp), 100 * C_CLK_PERIOD, 102 * C_CLK_PERIOD, ERROR, "2nd read should be executed 100 cycles after the first");

        log("\rFetch the 3rd result");
        await_completion(SBI_VVCT,2, v_cmd_idx+3, 2 * C_CLK_PERIOD, "3rd read should be executed 1 cycle after the 2nd");
        fetch_result(SBI_VVCT,2, v_cmd_idx+3, v_data, v_is_ok, "Fetching 3rd read-result");
        check_value(v_is_ok, ERROR, "Readback OK via fetch_result()");
        check_value(v_data(7 downto 0), x"C2", ERROR, "Readback data via fetch_result()");

        await_completion(SBI_VVCT, 2, 1000 ns);

      elsif run("read_of_executor_status_and_inter_bfm_delay") then
        log(ID_LOG_HDR, "Test of reading executor status");

        log("current_cmd_idx: " & to_string(shared_sbi_vvc_status(1).current_cmd_idx));
        log("previous_cmd_idx: " & to_string(shared_sbi_vvc_status(1).previous_cmd_idx));
        log("pending_cmd_cnt: " & to_string(shared_sbi_vvc_status(1).pending_cmd_cnt));
        check_value(shared_sbi_vvc_status(1).pending_cmd_cnt, 0, ERROR, "Checking that no commands are pending");
        sbi_write(SBI_VVCT,1, x"00", x"A0", "Write SBI1");
        sbi_write(SBI_VVCT,1, x"00", x"A0", "Write SBI1");
        sbi_write(SBI_VVCT,1, x"00", x"A0", "Write SBI1");
        log("current_cmd_idx: " & to_string(shared_sbi_vvc_status(1).current_cmd_idx));
        log("previous_cmd_idx: " & to_string(shared_sbi_vvc_status(1).previous_cmd_idx));
        check_value(shared_sbi_vvc_status(1).pending_cmd_cnt, 2, ERROR, "Checking pending commands");
        await_completion(SBI_VVCT,1,100 ns);
        log("current_cmd_idx: " & to_string(shared_sbi_vvc_status(1).current_cmd_idx));
        log("previous_cmd_idx: " & to_string(shared_sbi_vvc_status(1).previous_cmd_idx));
        check_value(shared_sbi_vvc_status(1).pending_cmd_cnt, 0, ERROR, "Checking that no commands are pending after completion");
        -- Cleanup
        sbi_write(SBI_VVCT,1, C_ADDR_FIFO_FLUSH, C_DATA_DONTCARE, "Flush FIFO 1");
        await_completion(SBI_VVCT,1,100 ns);

        log(ID_LOG_HDR, "Testing inter-bfm delay");

        log("\rChecking TIME_START2START");
        wait for C_CLK_PERIOD * 51;
        shared_sbi_vvc_config(1).inter_bfm_delay.delay_type := TIME_START2START;
        shared_sbi_vvc_config(1).inter_bfm_delay.delay_in_time := C_CLK_PERIOD * 50;
        v_timestamp := now;
        sbi_write(SBI_VVCT,1, x"00", x"A0", "First write to SBI1");
        sbi_write(SBI_VVCT,1, x"00", x"03", "Second write to SBI1");
        await_completion(SBI_VVCT, 1, 52 * C_CLK_PERIOD);
        check_value(((now - v_timestamp) = C_CLK_PERIOD*51), ERROR, "Checking that inter-bfm delay was upheld");

        log("\rChecking that insert_delay does not affect inter-BFM delay");
        wait for C_CLK_PERIOD * 51;
        v_timestamp := now;
        sbi_write(SBI_VVCT,1, x"00", x"AB", "First Write SBI1");
        insert_delay(SBI_VVCT,1, C_CLK_PERIOD);
        insert_delay(SBI_VVCT,1, C_CLK_PERIOD);
        insert_delay(SBI_VVCT,1, C_CLK_PERIOD);
        insert_delay(SBI_VVCT,1, C_CLK_PERIOD);
        sbi_write(SBI_VVCT,1, x"00", x"FF", "Second Write SBI1");
        await_completion(SBI_VVCT, 1, 52 * C_CLK_PERIOD + (4*C_CLK_PERIOD));
        check_value(((now - v_timestamp) = C_CLK_PERIOD*51 + (4*C_CLK_PERIOD)), ERROR, "Checking that inter-bfm delay was upheld");


        log("\rChecking TIME_FINISH2START");
        wait for C_CLK_PERIOD * 101;
        shared_sbi_vvc_config(1).inter_bfm_delay.delay_type := TIME_FINISH2START;
        shared_sbi_vvc_config(1).inter_bfm_delay.delay_in_time := C_CLK_PERIOD * 100;
        v_timestamp := now;
        sbi_write(SBI_VVCT,1, x"00", x"A0", "Write SBI1");
        sbi_write(SBI_VVCT,1, x"00", x"CC", "Write SBI1");
        await_completion(SBI_VVCT, 1, 103 * C_CLK_PERIOD);
        check_value(((now - v_timestamp) = C_CLK_PERIOD*102), ERROR, "Checking that inter-bfm delay was upheld");

        log("\rChecking TIME_START2START and provoking inter-bfm delay violation");
        wait for C_CLK_PERIOD * 10;
        increment_expected_alerts(TB_WARNING,2);
        shared_sbi_vvc_config(1).inter_bfm_delay.inter_bfm_delay_violation_severity := TB_WARNING;
        shared_sbi_vvc_config(1).inter_bfm_delay.delay_type := TIME_START2START;
        shared_sbi_vvc_config(1).inter_bfm_delay.delay_in_time := 1 ns;
        sbi_write(SBI_VVCT,1, x"00", x"A0", "First write to SBI1");
        sbi_write(SBI_VVCT,1, x"00", x"03", "Second write to SBI1");
        await_completion(SBI_VVCT, 1, 3 * C_CLK_PERIOD);

        log("Setting delay back to initial value");
        shared_sbi_vvc_config(1).inter_bfm_delay.delay_type := NO_DELAY;
        shared_sbi_vvc_config(1).inter_bfm_delay.delay_in_time := 0 ns;
        shared_sbi_vvc_config(1).inter_bfm_delay.inter_bfm_delay_violation_severity := WARNING;

      elsif run("distribution_of_vvc_commands") then
        log(ID_LOG_HDR, "Check that commands are distributed to the correct VVC channel");
        -- Calling an invalid channel will yield a TB_WARNING from each of the UART channels
        -- We will also get another TB_WARNING from the timeout, related to having more decimals in the log time than we can display
        increment_expected_alerts(TB_WARNING,3);
        -- Calling an invalid channel will also cause a timeout, since the target VVC does not exist. This results in an ERROR
        increment_expected_alerts(TB_ERROR,3);
        insert_delay(SBI_VVCT, 1, TX, C_CLK_PERIOD, "Inserting delay on SBI TX channel, expecting tb warning and tb error");
        insert_delay(SBI_VVCT, 1, RX, C_CLK_PERIOD, "Inserting delay on SBI RX channel, expecting tb warning and tb error");
        insert_delay(SBI_VVCT, 42, C_CLK_PERIOD, "Inserting delay on SBI VVC 42, expecting tb error");
        log("Logging a message to provoke the tb warning due to truncated timestamp");

      elsif run("vvc_broadcast_test") then
        log(ID_LOG_HDR, "Check that commands are distributed to the correct VVC channel");

        enable_log_msg(VVC_BROADCAST, ALL_MESSAGES);

        -- Fill FIFO 1
        sbi_write(SBI_VVCT,C_VVCT_ALL_INSTANCES, C_ADDR_FIFO_PUT, x"01", "Write PUT on both FIFOs");
        sbi_write(SBI_VVCT,C_VVCT_ALL_INSTANCES, C_ADDR_FIFO_PUT, x"56", "Write PUT on both FIFOs");
        sbi_write(SBI_VVCT,C_VVCT_ALL_INSTANCES, C_ADDR_FIFO_PUT, x"a3", "Write PUT on both FIFOs");
        sbi_write(SBI_VVCT,C_VVCT_ALL_INSTANCES, C_ADDR_FIFO_PUT, x"4d", "Write PUT on both FIFOs");
        sbi_write(SBI_VVCT,C_VVCT_ALL_INSTANCES, C_ADDR_FIFO_PUT, x"00", "Write PUT on both FIFOs");
        sbi_write(SBI_VVCT,C_VVCT_ALL_INSTANCES, C_ADDR_FIFO_PUT, x"42", "Write PUT on both FIFOs");
        await_completion(SBI_VVCT,C_VVCT_ALL_INSTANCES, 1000 ns, "Await execution for both VVCs");

        -- Poll from FIFO 1
        sbi_poll_until(SBI_VVCT,1, C_ADDR_FIFO_GET,  x"42", "Test of POLL_UNTIL within 100 ns", 0, 100 ns, ERROR);

        -- Poll from FIFO 2
        sbi_poll_until(SBI_VVCT,2, C_ADDR_FIFO_GET,  x"42", "Test of POLL_UNTIL within 10 occurrences", 10, 0 ns, ERROR);

        await_completion(SBI_VVCT,C_VVCT_ALL_INSTANCES, 1000 ns, "Await execution");

        log(ID_LOG_HDR, "Checking broadcast of flush_command_queue");
        sbi_write(SBI_VVCT,C_VVCT_ALL_INSTANCES, C_ADDR_FIFO_PUT, x"4d", "Write PUT on both FIFOs");
        sbi_write(SBI_VVCT,C_VVCT_ALL_INSTANCES, C_ADDR_FIFO_PUT, x"00", "Write PUT on both FIFOs");
        sbi_write(SBI_VVCT,C_VVCT_ALL_INSTANCES, C_ADDR_FIFO_PUT, x"42", "Write PUT on both FIFOs");
        flush_command_queue(VVC_BROADCAST, "Flushing all commands");
        await_completion(SBI_VVCT,C_VVCT_ALL_INSTANCES, 2*C_CLK_PERIOD, "Await flush completion");


        log(ID_LOG_HDR, "Checking broadcast of insert_delay (time)");

        log("Setting no initial inter-bfm delay");
        shared_sbi_vvc_config(1).inter_bfm_delay.delay_type := NO_DELAY;
        shared_sbi_vvc_config(1).inter_bfm_delay.delay_in_time := 0 ns;
        shared_sbi_vvc_config(1).inter_bfm_delay.inter_bfm_delay_violation_severity := WARNING;

        v_timestamp := now;
        sbi_write(SBI_VVCT,C_VVCT_ALL_INSTANCES, x"00", x"AB", "First Write SBI1");
        insert_delay(VVC_BROADCAST, C_CLK_PERIOD, "Inserting delay in all VVCs");
        insert_delay(VVC_BROADCAST, C_CLK_PERIOD, "Inserting delay in all VVCs");
        insert_delay(VVC_BROADCAST, C_CLK_PERIOD, "Inserting delay in all VVCs");
        insert_delay(VVC_BROADCAST, C_CLK_PERIOD, "Inserting delay in all VVCs");
        sbi_write(SBI_VVCT,C_VVCT_ALL_INSTANCES, x"00", x"FF", "Second Write SBI1");
        await_completion(SBI_VVCT, 1, 7 * C_CLK_PERIOD);
        check_value(((now - v_timestamp) = C_CLK_PERIOD*6), ERROR, "Checking that inter-bfm delay was upheld");

        await_completion(SBI_VVCT,2, 1000 ns, "Await execution");

      elsif run("vvc_setup_and_hold_time_test") then
        log(ID_LOG_HDR, "Checking setup and hold time");

        -- Set setup and hold times
        log("Setup time: 2 ns, hold time: 1 ns");
        shared_sbi_vvc_config(1).bfm_config.setup_time := 2 ns;
        shared_sbi_vvc_config(1).bfm_config.hold_time := 1 ns;

        -- Check for sbi_write
        sbi_write(SBI_VVCT,1, x"00", x"AA", "Write SBI1");
        await_value(sbi1_if.wena, '1', 0 ns, 100 ns, ERROR, "Waiting on wena from SBI1");
        await_value(clk, '1', 2 ns, 2.01 ns, ERROR, "Waiting on positive clk edge, shall occour 2 ns after wdata");
        check_value(sbi1_if.wena'last_event, 2 ns, ERROR, "Check setup time", C_SCOPE, ID_SEQUENCER);
        await_value(sbi1_if.wena, '0', 1 ns, 1.01 ns, ERROR, "Waiting on wena to go inactive, should occuer after 1 ns");
        check_value(clk'last_event, 1 ns, ERROR, "Check hold time", C_SCOPE, ID_SEQUENCER);

        -- Check for sbi_read
        sbi_read(SBI_VVCT,1, C_ADDR_FIFO_COUNT, "Readback inside VVC");
        await_value(sbi1_if.rena, '1', 0 ns, 100 ns, ERROR, "Waiting on rena from SBI1");
        await_value(clk, '1', 2 ns, 2.01 ns, ERROR, "Waiting on positive clk edge, shall occour 2 ns after wdata");
        check_value(sbi1_if.rena'last_event, 2 ns, ERROR, "Check setup time", C_SCOPE, ID_SEQUENCER);
        await_value(sbi1_if.rena, '0', 1 ns, 1.01 ns, ERROR, "Waiting on rena to go inactive, should occuer after 1 ns");
        check_value(clk'last_event, 1 ns, ERROR, "Check hold time", C_SCOPE, ID_SEQUENCER);

        -- New values
        -- Set setup and hold times
        log("\nSetup time: 1 ns, hold time: 3 ns");
        shared_sbi_vvc_config(1).bfm_config.setup_time := 1 ns;
        shared_sbi_vvc_config(1).bfm_config.hold_time := 3 ns;

        -- Check for sbi_write
        sbi_write(SBI_VVCT,1, x"00", x"AB", "Write SBI1");
        await_value(sbi1_if.wena, '1', 0 ns, 100 ns, ERROR, "Waiting on wena from SBI1");
        await_value(clk, '1', 1 ns, 1.01 ns, ERROR, "Waiting on positive clk edge, shall occour 1 ns after wdata");
        check_value(sbi1_if.wena'last_event, 1 ns, ERROR, "Check setup time", C_SCOPE, ID_SEQUENCER);
        await_value(sbi1_if.wena, '0', 3 ns, 3.01 ns, ERROR, "Waiting on wena to go inactive, should occuer after 3 ns");
        check_value(clk'last_event, 3 ns, ERROR, "Check hold time", C_SCOPE, ID_SEQUENCER);

        -- Check for sbi_read
        sbi_read(SBI_VVCT,1, C_ADDR_FIFO_COUNT, "Readback inside VVC");
        await_value(sbi1_if.rena, '1', 0 ns, 100 ns, ERROR, "Waiting on rena from SBI1");
        await_value(clk, '1', 1 ns, 1.01 ns, ERROR, "Waiting on positive clk edge, shall occour 2 ns after wdata");
        check_value(sbi1_if.rena'last_event, 1 ns, ERROR, "Check setup time", C_SCOPE, ID_SEQUENCER);
        await_value(sbi1_if.rena, '0', 3 ns, 3.01 ns, ERROR, "Waiting on rena to go inactive, should occuer after 1 ns");
        check_value(clk'last_event, 3 ns, ERROR, "Check hold time", C_SCOPE, ID_SEQUENCER);

      end if;
    end loop;
    --==================================================================================================
    -- Ending the simulation
    --------------------------------------------------------------------------------------
    wait for 1000 ns;  -- to allow some time for completion
    report_alert_counters(VOID);
    log(ID_LOG_HDR, "SIMULATION COMPLETED");

    -- Cleanup VUnit. The UVVM-Util error status is imported into VUnit at this
    -- point. This is neccessary when the UVVM-Util alert stop limit is set such that
    -- UVVM-Util doesn't stop on the first error. In that case VUnit has no way of
    -- knowing the error status unless you tell it.
    for alert_level in NOTE to t_alert_level'right loop
      if alert_level /= MANUAL_CHECK and get_alert_counter(alert_level, REGARD) /= get_alert_counter(alert_level, EXPECT) then
        v_alert_num_mismatch := true;
      end if;
    end loop;

    test_runner_cleanup(runner, v_alert_num_mismatch);
    wait;

  end process p_main;

end func;
