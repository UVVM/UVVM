-------------------------------------------------------
--  Copyright (c) 1995/2006 Xilinx Inc.
--  All Right Reserved.
-------------------------------------------------------
--
--   ____  ____
--  /   /\/   / 
-- /___/  \  /     Vendor      : Xilinx 
-- \   \   \/      Version : 11.1
--  \   \          Description : 
--  /   /                      
-- /___/   /\      Filename    : PPC440.vhd
-- \   \  /  \     Timestamp   : Thu Apr 19 15:56:12 2007

--  \__ \/\__ \                   
--                                 
--  Generated by    : write_vhdl
--  Revision: 
-------------------------------------------------------

----- CELL PPC440 -----

library IEEE;
use IEEE.STD_LOGIC_1164.all;

library IEEE;
use IEEE.VITAL_Timing.all;

library unisim;
use unisim.VCOMPONENTS.all;

library secureip;
use secureip.all;

entity PPC440 is
generic (
	APU_CONTROL : bit_vector := X"02000";
	APU_UDI0 : bit_vector := X"000000";
	APU_UDI1 : bit_vector := X"000000";
	APU_UDI10 : bit_vector := X"000000";
	APU_UDI11 : bit_vector := X"000000";
	APU_UDI12 : bit_vector := X"000000";
	APU_UDI13 : bit_vector := X"000000";
	APU_UDI14 : bit_vector := X"000000";
	APU_UDI15 : bit_vector := X"000000";
	APU_UDI2 : bit_vector := X"000000";
	APU_UDI3 : bit_vector := X"000000";
	APU_UDI4 : bit_vector := X"000000";
	APU_UDI5 : bit_vector := X"000000";
	APU_UDI6 : bit_vector := X"000000";
	APU_UDI7 : bit_vector := X"000000";
	APU_UDI8 : bit_vector := X"000000";
	APU_UDI9 : bit_vector := X"000000";
	CLOCK_DELAY : boolean := FALSE;
	DCR_AUTOLOCK_ENABLE : boolean := TRUE;
	DMA0_CONTROL : bit_vector := X"00";
	DMA0_RXCHANNELCTRL : bit_vector := X"01010000";
	DMA0_RXIRQTIMER : bit_vector := X"3FF";
	DMA0_TXCHANNELCTRL : bit_vector := X"01010000";
	DMA0_TXIRQTIMER : bit_vector := X"3FF";
	DMA1_CONTROL : bit_vector := X"00";
	DMA1_RXCHANNELCTRL : bit_vector := X"01010000";
	DMA1_RXIRQTIMER : bit_vector := X"3FF";
	DMA1_TXCHANNELCTRL : bit_vector := X"01010000";
	DMA1_TXIRQTIMER : bit_vector := X"3FF";
	DMA2_CONTROL : bit_vector := X"00";
	DMA2_RXCHANNELCTRL : bit_vector := X"01010000";
	DMA2_RXIRQTIMER : bit_vector := X"3FF";
	DMA2_TXCHANNELCTRL : bit_vector := X"01010000";
	DMA2_TXIRQTIMER : bit_vector := X"3FF";
	DMA3_CONTROL : bit_vector := X"00";
	DMA3_RXCHANNELCTRL : bit_vector := X"01010000";
	DMA3_RXIRQTIMER : bit_vector := X"3FF";
	DMA3_TXCHANNELCTRL : bit_vector := X"01010000";
	DMA3_TXIRQTIMER : bit_vector := X"3FF";
	INTERCONNECT_IMASK : bit_vector := X"FFFFFFFF";
	INTERCONNECT_TMPL_SEL : bit_vector := X"3FFFFFFF";
	MI_ARBCONFIG : bit_vector := X"00432010";
	MI_BANKCONFLICT_MASK : bit_vector := X"00000000";
	MI_CONTROL : bit_vector := X"0000008F";
	MI_ROWCONFLICT_MASK : bit_vector := X"00000000";
	PPCDM_ASYNCMODE : boolean := FALSE;
	PPCDS_ASYNCMODE : boolean := FALSE;
	PPCM_ARBCONFIG : bit_vector := X"00432010";
	PPCM_CONTROL : bit_vector := X"8000009F";
	PPCM_COUNTER : bit_vector := X"00000500";
	PPCS0_ADDRMAP_TMPL0 : bit_vector := X"FFFFFFFF";
	PPCS0_ADDRMAP_TMPL1 : bit_vector := X"FFFFFFFF";
	PPCS0_ADDRMAP_TMPL2 : bit_vector := X"FFFFFFFF";
	PPCS0_ADDRMAP_TMPL3 : bit_vector := X"FFFFFFFF";
	PPCS0_CONTROL : bit_vector := X"8033336C";
	PPCS0_WIDTH_128N64 : boolean := TRUE;
	PPCS1_ADDRMAP_TMPL0 : bit_vector := X"FFFFFFFF";
	PPCS1_ADDRMAP_TMPL1 : bit_vector := X"FFFFFFFF";
	PPCS1_ADDRMAP_TMPL2 : bit_vector := X"FFFFFFFF";
	PPCS1_ADDRMAP_TMPL3 : bit_vector := X"FFFFFFFF";
	PPCS1_CONTROL : bit_vector := X"8033336C";
	PPCS1_WIDTH_128N64 : boolean := TRUE;
	XBAR_ADDRMAP_TMPL0 : bit_vector := X"FFFF0000";
	XBAR_ADDRMAP_TMPL1 : bit_vector := X"00000000";
	XBAR_ADDRMAP_TMPL2 : bit_vector := X"00000000";
	XBAR_ADDRMAP_TMPL3 : bit_vector := X"00000000"




  );

port (
		APUFCMDECFPUOP : out std_ulogic;
		APUFCMDECLDSTXFERSIZE : out std_logic_vector(0 to 2);
		APUFCMDECLOAD : out std_ulogic;
		APUFCMDECNONAUTON : out std_ulogic;
		APUFCMDECSTORE : out std_ulogic;
		APUFCMDECUDI : out std_logic_vector(0 to 3);
		APUFCMDECUDIVALID : out std_ulogic;
		APUFCMENDIAN : out std_ulogic;
		APUFCMFLUSH : out std_ulogic;
		APUFCMINSTRUCTION : out std_logic_vector(0 to 31);
		APUFCMINSTRVALID : out std_ulogic;
		APUFCMLOADBYTEADDR : out std_logic_vector(0 to 3);
		APUFCMLOADDATA : out std_logic_vector(0 to 127);
		APUFCMLOADDVALID : out std_ulogic;
		APUFCMMSRFE0 : out std_ulogic;
		APUFCMMSRFE1 : out std_ulogic;
		APUFCMNEXTINSTRREADY : out std_ulogic;
		APUFCMOPERANDVALID : out std_ulogic;
		APUFCMRADATA : out std_logic_vector(0 to 31);
		APUFCMRBDATA : out std_logic_vector(0 to 31);
		APUFCMWRITEBACKOK : out std_ulogic;
		C440CPMCORESLEEPREQ : out std_ulogic;
		C440CPMDECIRPTREQ : out std_ulogic;
		C440CPMFITIRPTREQ : out std_ulogic;
		C440CPMMSRCE : out std_ulogic;
		C440CPMMSREE : out std_ulogic;
		C440CPMTIMERRESETREQ : out std_ulogic;
		C440CPMWDIRPTREQ : out std_ulogic;
		C440DBGSYSTEMCONTROL : out std_logic_vector(0 to 7);
		C440JTGTDO : out std_ulogic;
		C440JTGTDOEN : out std_ulogic;
		C440MACHINECHECK : out std_ulogic;
		C440RSTCHIPRESETREQ : out std_ulogic;
		C440RSTCORERESETREQ : out std_ulogic;
		C440RSTSYSTEMRESETREQ : out std_ulogic;
		C440TRCBRANCHSTATUS : out std_logic_vector(0 to 2);
		C440TRCCYCLE : out std_ulogic;
		C440TRCEXECUTIONSTATUS : out std_logic_vector(0 to 4);
		C440TRCTRACESTATUS : out std_logic_vector(0 to 6);
		C440TRCTRIGGEREVENTOUT : out std_ulogic;
		C440TRCTRIGGEREVENTTYPE : out std_logic_vector(0 to 13);
		DMA0LLRSTENGINEACK : out std_ulogic;
		DMA0LLRXDSTRDYN : out std_ulogic;
		DMA0LLTXD : out std_logic_vector(0 to 31);
		DMA0LLTXEOFN : out std_ulogic;
		DMA0LLTXEOPN : out std_ulogic;
		DMA0LLTXREM : out std_logic_vector(0 to 3);
		DMA0LLTXSOFN : out std_ulogic;
		DMA0LLTXSOPN : out std_ulogic;
		DMA0LLTXSRCRDYN : out std_ulogic;
		DMA0RXIRQ : out std_ulogic;
		DMA0TXIRQ : out std_ulogic;
		DMA1LLRSTENGINEACK : out std_ulogic;
		DMA1LLRXDSTRDYN : out std_ulogic;
		DMA1LLTXD : out std_logic_vector(0 to 31);
		DMA1LLTXEOFN : out std_ulogic;
		DMA1LLTXEOPN : out std_ulogic;
		DMA1LLTXREM : out std_logic_vector(0 to 3);
		DMA1LLTXSOFN : out std_ulogic;
		DMA1LLTXSOPN : out std_ulogic;
		DMA1LLTXSRCRDYN : out std_ulogic;
		DMA1RXIRQ : out std_ulogic;
		DMA1TXIRQ : out std_ulogic;
		DMA2LLRSTENGINEACK : out std_ulogic;
		DMA2LLRXDSTRDYN : out std_ulogic;
		DMA2LLTXD : out std_logic_vector(0 to 31);
		DMA2LLTXEOFN : out std_ulogic;
		DMA2LLTXEOPN : out std_ulogic;
		DMA2LLTXREM : out std_logic_vector(0 to 3);
		DMA2LLTXSOFN : out std_ulogic;
		DMA2LLTXSOPN : out std_ulogic;
		DMA2LLTXSRCRDYN : out std_ulogic;
		DMA2RXIRQ : out std_ulogic;
		DMA2TXIRQ : out std_ulogic;
		DMA3LLRSTENGINEACK : out std_ulogic;
		DMA3LLRXDSTRDYN : out std_ulogic;
		DMA3LLTXD : out std_logic_vector(0 to 31);
		DMA3LLTXEOFN : out std_ulogic;
		DMA3LLTXEOPN : out std_ulogic;
		DMA3LLTXREM : out std_logic_vector(0 to 3);
		DMA3LLTXSOFN : out std_ulogic;
		DMA3LLTXSOPN : out std_ulogic;
		DMA3LLTXSRCRDYN : out std_ulogic;
		DMA3RXIRQ : out std_ulogic;
		DMA3TXIRQ : out std_ulogic;
		MIMCADDRESS : out std_logic_vector(0 to 35);
		MIMCADDRESSVALID : out std_ulogic;
		MIMCBANKCONFLICT : out std_ulogic;
		MIMCBYTEENABLE : out std_logic_vector(0 to 15);
		MIMCREADNOTWRITE : out std_ulogic;
		MIMCROWCONFLICT : out std_ulogic;
		MIMCWRITEDATA : out std_logic_vector(0 to 127);
		MIMCWRITEDATAVALID : out std_ulogic;
		PPCCPMINTERCONNECTBUSY : out std_ulogic;
		PPCDMDCRABUS : out std_logic_vector(0 to 9);
		PPCDMDCRDBUSOUT : out std_logic_vector(0 to 31);
		PPCDMDCRREAD : out std_ulogic;
		PPCDMDCRUABUS : out std_logic_vector(20 to 21);
		PPCDMDCRWRITE : out std_ulogic;
		PPCDSDCRACK : out std_ulogic;
		PPCDSDCRDBUSIN : out std_logic_vector(0 to 31);
		PPCDSDCRTIMEOUTWAIT : out std_ulogic;
		PPCEICINTERCONNECTIRQ : out std_ulogic;
		PPCMPLBABORT : out std_ulogic;
		PPCMPLBABUS : out std_logic_vector(0 to 31);
		PPCMPLBBE : out std_logic_vector(0 to 15);
		PPCMPLBBUSLOCK : out std_ulogic;
		PPCMPLBLOCKERR : out std_ulogic;
		PPCMPLBPRIORITY : out std_logic_vector(0 to 1);
		PPCMPLBRDBURST : out std_ulogic;
		PPCMPLBREQUEST : out std_ulogic;
		PPCMPLBRNW : out std_ulogic;
		PPCMPLBSIZE : out std_logic_vector(0 to 3);
		PPCMPLBTATTRIBUTE : out std_logic_vector(0 to 15);
		PPCMPLBTYPE : out std_logic_vector(0 to 2);
		PPCMPLBUABUS : out std_logic_vector(28 to 31);
		PPCMPLBWRBURST : out std_ulogic;
		PPCMPLBWRDBUS : out std_logic_vector(0 to 127);
		PPCS0PLBADDRACK : out std_ulogic;
		PPCS0PLBMBUSY : out std_logic_vector(0 to 3);
		PPCS0PLBMIRQ : out std_logic_vector(0 to 3);
		PPCS0PLBMRDERR : out std_logic_vector(0 to 3);
		PPCS0PLBMWRERR : out std_logic_vector(0 to 3);
		PPCS0PLBRDBTERM : out std_ulogic;
		PPCS0PLBRDCOMP : out std_ulogic;
		PPCS0PLBRDDACK : out std_ulogic;
		PPCS0PLBRDDBUS : out std_logic_vector(0 to 127);
		PPCS0PLBRDWDADDR : out std_logic_vector(0 to 3);
		PPCS0PLBREARBITRATE : out std_ulogic;
		PPCS0PLBSSIZE : out std_logic_vector(0 to 1);
		PPCS0PLBWAIT : out std_ulogic;
		PPCS0PLBWRBTERM : out std_ulogic;
		PPCS0PLBWRCOMP : out std_ulogic;
		PPCS0PLBWRDACK : out std_ulogic;
		PPCS1PLBADDRACK : out std_ulogic;
		PPCS1PLBMBUSY : out std_logic_vector(0 to 3);
		PPCS1PLBMIRQ : out std_logic_vector(0 to 3);
		PPCS1PLBMRDERR : out std_logic_vector(0 to 3);
		PPCS1PLBMWRERR : out std_logic_vector(0 to 3);
		PPCS1PLBRDBTERM : out std_ulogic;
		PPCS1PLBRDCOMP : out std_ulogic;
		PPCS1PLBRDDACK : out std_ulogic;
		PPCS1PLBRDDBUS : out std_logic_vector(0 to 127);
		PPCS1PLBRDWDADDR : out std_logic_vector(0 to 3);
		PPCS1PLBREARBITRATE : out std_ulogic;
		PPCS1PLBSSIZE : out std_logic_vector(0 to 1);
		PPCS1PLBWAIT : out std_ulogic;
		PPCS1PLBWRBTERM : out std_ulogic;
		PPCS1PLBWRCOMP : out std_ulogic;
		PPCS1PLBWRDACK : out std_ulogic;

		CPMC440CLK : in std_ulogic;
		CPMC440CLKEN : in std_ulogic;
		CPMC440CORECLOCKINACTIVE : in std_ulogic;
		CPMC440TIMERCLOCK : in std_ulogic;
		CPMDCRCLK : in std_ulogic;
		CPMDMA0LLCLK : in std_ulogic;
		CPMDMA1LLCLK : in std_ulogic;
		CPMDMA2LLCLK : in std_ulogic;
		CPMDMA3LLCLK : in std_ulogic;
		CPMFCMCLK : in std_ulogic;
		CPMINTERCONNECTCLK : in std_ulogic;
		CPMINTERCONNECTCLKEN : in std_ulogic;
		CPMINTERCONNECTCLKNTO1 : in std_ulogic;
		CPMMCCLK : in std_ulogic;
		CPMPPCMPLBCLK : in std_ulogic;
		CPMPPCS0PLBCLK : in std_ulogic;
		CPMPPCS1PLBCLK : in std_ulogic;
		DBGC440DEBUGHALT : in std_ulogic;
		DBGC440SYSTEMSTATUS : in std_logic_vector(0 to 4);
		DBGC440UNCONDDEBUGEVENT : in std_ulogic;
		DCRPPCDMACK : in std_ulogic;
		DCRPPCDMDBUSIN : in std_logic_vector(0 to 31);
		DCRPPCDMTIMEOUTWAIT : in std_ulogic;
		DCRPPCDSABUS : in std_logic_vector(0 to 9);
		DCRPPCDSDBUSOUT : in std_logic_vector(0 to 31);
		DCRPPCDSREAD : in std_ulogic;
		DCRPPCDSWRITE : in std_ulogic;
		EICC440CRITIRQ : in std_ulogic;
		EICC440EXTIRQ : in std_ulogic;
		FCMAPUCONFIRMINSTR : in std_ulogic;
		FCMAPUCR : in std_logic_vector(0 to 3);
		FCMAPUDONE : in std_ulogic;
		FCMAPUEXCEPTION : in std_ulogic;
		FCMAPUFPSCRFEX : in std_ulogic;
		FCMAPURESULT : in std_logic_vector(0 to 31);
		FCMAPURESULTVALID : in std_ulogic;
		FCMAPUSLEEPNOTREADY : in std_ulogic;
		FCMAPUSTOREDATA : in std_logic_vector(0 to 127);
		JTGC440TCK : in std_ulogic;
		JTGC440TDI : in std_ulogic;
		JTGC440TMS : in std_ulogic;
		JTGC440TRSTNEG : in std_ulogic;
		LLDMA0RSTENGINEREQ : in std_ulogic;
		LLDMA0RXD : in std_logic_vector(0 to 31);
		LLDMA0RXEOFN : in std_ulogic;
		LLDMA0RXEOPN : in std_ulogic;
		LLDMA0RXREM : in std_logic_vector(0 to 3);
		LLDMA0RXSOFN : in std_ulogic;
		LLDMA0RXSOPN : in std_ulogic;
		LLDMA0RXSRCRDYN : in std_ulogic;
		LLDMA0TXDSTRDYN : in std_ulogic;
		LLDMA1RSTENGINEREQ : in std_ulogic;
		LLDMA1RXD : in std_logic_vector(0 to 31);
		LLDMA1RXEOFN : in std_ulogic;
		LLDMA1RXEOPN : in std_ulogic;
		LLDMA1RXREM : in std_logic_vector(0 to 3);
		LLDMA1RXSOFN : in std_ulogic;
		LLDMA1RXSOPN : in std_ulogic;
		LLDMA1RXSRCRDYN : in std_ulogic;
		LLDMA1TXDSTRDYN : in std_ulogic;
		LLDMA2RSTENGINEREQ : in std_ulogic;
		LLDMA2RXD : in std_logic_vector(0 to 31);
		LLDMA2RXEOFN : in std_ulogic;
		LLDMA2RXEOPN : in std_ulogic;
		LLDMA2RXREM : in std_logic_vector(0 to 3);
		LLDMA2RXSOFN : in std_ulogic;
		LLDMA2RXSOPN : in std_ulogic;
		LLDMA2RXSRCRDYN : in std_ulogic;
		LLDMA2TXDSTRDYN : in std_ulogic;
		LLDMA3RSTENGINEREQ : in std_ulogic;
		LLDMA3RXD : in std_logic_vector(0 to 31);
		LLDMA3RXEOFN : in std_ulogic;
		LLDMA3RXEOPN : in std_ulogic;
		LLDMA3RXREM : in std_logic_vector(0 to 3);
		LLDMA3RXSOFN : in std_ulogic;
		LLDMA3RXSOPN : in std_ulogic;
		LLDMA3RXSRCRDYN : in std_ulogic;
		LLDMA3TXDSTRDYN : in std_ulogic;
		MCMIADDRREADYTOACCEPT : in std_ulogic;
		MCMIREADDATA : in std_logic_vector(0 to 127);
		MCMIREADDATAERR : in std_ulogic;
		MCMIREADDATAVALID : in std_ulogic;
		PLBPPCMADDRACK : in std_ulogic;
		PLBPPCMMBUSY : in std_ulogic;
		PLBPPCMMIRQ : in std_ulogic;
		PLBPPCMMRDERR : in std_ulogic;
		PLBPPCMMWRERR : in std_ulogic;
		PLBPPCMRDBTERM : in std_ulogic;
		PLBPPCMRDDACK : in std_ulogic;
		PLBPPCMRDDBUS : in std_logic_vector(0 to 127);
		PLBPPCMRDPENDPRI : in std_logic_vector(0 to 1);
		PLBPPCMRDPENDREQ : in std_ulogic;
		PLBPPCMRDWDADDR : in std_logic_vector(0 to 3);
		PLBPPCMREARBITRATE : in std_ulogic;
		PLBPPCMREQPRI : in std_logic_vector(0 to 1);
		PLBPPCMSSIZE : in std_logic_vector(0 to 1);
		PLBPPCMTIMEOUT : in std_ulogic;
		PLBPPCMWRBTERM : in std_ulogic;
		PLBPPCMWRDACK : in std_ulogic;
		PLBPPCMWRPENDPRI : in std_logic_vector(0 to 1);
		PLBPPCMWRPENDREQ : in std_ulogic;
		PLBPPCS0ABORT : in std_ulogic;
		PLBPPCS0ABUS : in std_logic_vector(0 to 31);
		PLBPPCS0BE : in std_logic_vector(0 to 15);
		PLBPPCS0BUSLOCK : in std_ulogic;
		PLBPPCS0LOCKERR : in std_ulogic;
		PLBPPCS0MASTERID : in std_logic_vector(0 to 1);
		PLBPPCS0MSIZE : in std_logic_vector(0 to 1);
		PLBPPCS0PAVALID : in std_ulogic;
		PLBPPCS0RDBURST : in std_ulogic;
		PLBPPCS0RDPENDPRI : in std_logic_vector(0 to 1);
		PLBPPCS0RDPENDREQ : in std_ulogic;
		PLBPPCS0RDPRIM : in std_ulogic;
		PLBPPCS0REQPRI : in std_logic_vector(0 to 1);
		PLBPPCS0RNW : in std_ulogic;
		PLBPPCS0SAVALID : in std_ulogic;
		PLBPPCS0SIZE : in std_logic_vector(0 to 3);
		PLBPPCS0TATTRIBUTE : in std_logic_vector(0 to 15);
		PLBPPCS0TYPE : in std_logic_vector(0 to 2);
		PLBPPCS0UABUS : in std_logic_vector(28 to 31);
		PLBPPCS0WRBURST : in std_ulogic;
		PLBPPCS0WRDBUS : in std_logic_vector(0 to 127);
		PLBPPCS0WRPENDPRI : in std_logic_vector(0 to 1);
		PLBPPCS0WRPENDREQ : in std_ulogic;
		PLBPPCS0WRPRIM : in std_ulogic;
		PLBPPCS1ABORT : in std_ulogic;
		PLBPPCS1ABUS : in std_logic_vector(0 to 31);
		PLBPPCS1BE : in std_logic_vector(0 to 15);
		PLBPPCS1BUSLOCK : in std_ulogic;
		PLBPPCS1LOCKERR : in std_ulogic;
		PLBPPCS1MASTERID : in std_logic_vector(0 to 1);
		PLBPPCS1MSIZE : in std_logic_vector(0 to 1);
		PLBPPCS1PAVALID : in std_ulogic;
		PLBPPCS1RDBURST : in std_ulogic;
		PLBPPCS1RDPENDPRI : in std_logic_vector(0 to 1);
		PLBPPCS1RDPENDREQ : in std_ulogic;
		PLBPPCS1RDPRIM : in std_ulogic;
		PLBPPCS1REQPRI : in std_logic_vector(0 to 1);
		PLBPPCS1RNW : in std_ulogic;
		PLBPPCS1SAVALID : in std_ulogic;
		PLBPPCS1SIZE : in std_logic_vector(0 to 3);
		PLBPPCS1TATTRIBUTE : in std_logic_vector(0 to 15);
		PLBPPCS1TYPE : in std_logic_vector(0 to 2);
		PLBPPCS1UABUS : in std_logic_vector(28 to 31);
		PLBPPCS1WRBURST : in std_ulogic;
		PLBPPCS1WRDBUS : in std_logic_vector(0 to 127);
		PLBPPCS1WRPENDPRI : in std_logic_vector(0 to 1);
		PLBPPCS1WRPENDREQ : in std_ulogic;
		PLBPPCS1WRPRIM : in std_ulogic;
		RSTC440RESETCHIP : in std_ulogic;
		RSTC440RESETCORE : in std_ulogic;
		RSTC440RESETSYSTEM : in std_ulogic;
		TIEC440DCURDLDCACHEPLBPRIO : in std_logic_vector(0 to 1);
		TIEC440DCURDNONCACHEPLBPRIO : in std_logic_vector(0 to 1);
		TIEC440DCURDTOUCHPLBPRIO : in std_logic_vector(0 to 1);
		TIEC440DCURDURGENTPLBPRIO : in std_logic_vector(0 to 1);
		TIEC440DCUWRFLUSHPLBPRIO : in std_logic_vector(0 to 1);
		TIEC440DCUWRSTOREPLBPRIO : in std_logic_vector(0 to 1);
		TIEC440DCUWRURGENTPLBPRIO : in std_logic_vector(0 to 1);
		TIEC440ENDIANRESET : in std_ulogic;
		TIEC440ERPNRESET : in std_logic_vector(0 to 3);
		TIEC440ICURDFETCHPLBPRIO : in std_logic_vector(0 to 1);
		TIEC440ICURDSPECPLBPRIO : in std_logic_vector(0 to 1);
		TIEC440ICURDTOUCHPLBPRIO : in std_logic_vector(0 to 1);
		TIEC440PIR : in std_logic_vector(28 to 31);
		TIEC440PVR : in std_logic_vector(28 to 31);
		TIEC440USERRESET : in std_logic_vector(0 to 3);
		TIEDCRBASEADDR : in std_logic_vector(0 to 1);
		TRCC440TRACEDISABLE : in std_ulogic;
		TRCC440TRIGGEREVENTIN : in std_ulogic
     );
end PPC440;

architecture PPC440_V of PPC440 is

  component PPC440_SWIFT
    port (
      APUFCMDECFPUOP       : out std_ulogic;
      APUFCMDECLDSTXFERSIZE : out std_logic_vector(0 to 2);
      APUFCMDECLOAD        : out std_ulogic;
      APUFCMDECNONAUTON    : out std_ulogic;
      APUFCMDECSTORE       : out std_ulogic;
      APUFCMDECUDI         : out std_logic_vector(0 to 3);
      APUFCMDECUDIVALID    : out std_ulogic;
      APUFCMENDIAN         : out std_ulogic;
      APUFCMFLUSH          : out std_ulogic;
      APUFCMINSTRUCTION    : out std_logic_vector(0 to 31);
      APUFCMINSTRVALID     : out std_ulogic;
      APUFCMLOADBYTEADDR   : out std_logic_vector(0 to 3);
      APUFCMLOADDATA       : out std_logic_vector(0 to 127);
      APUFCMLOADDVALID     : out std_ulogic;
      APUFCMMSRFE0         : out std_ulogic;
      APUFCMMSRFE1         : out std_ulogic;
      APUFCMNEXTINSTRREADY : out std_ulogic;
      APUFCMOPERANDVALID   : out std_ulogic;
      APUFCMRADATA         : out std_logic_vector(0 to 31);
      APUFCMRBDATA         : out std_logic_vector(0 to 31);
      APUFCMWRITEBACKOK    : out std_ulogic;
      C440CPMCORESLEEPREQ  : out std_ulogic;
      C440CPMDECIRPTREQ    : out std_ulogic;
      C440CPMFITIRPTREQ    : out std_ulogic;
      C440CPMMSRCE         : out std_ulogic;
      C440CPMMSREE         : out std_ulogic;
      C440CPMTIMERRESETREQ : out std_ulogic;
      C440CPMWDIRPTREQ     : out std_ulogic;
      C440DBGSYSTEMCONTROL : out std_logic_vector(0 to 7);
      C440JTGTDO           : out std_ulogic;
      C440JTGTDOEN         : out std_ulogic;
      C440MACHINECHECK     : out std_ulogic;
      C440RSTCHIPRESETREQ  : out std_ulogic;
      C440RSTCORERESETREQ  : out std_ulogic;
      C440RSTSYSTEMRESETREQ : out std_ulogic;
      C440TRCBRANCHSTATUS  : out std_logic_vector(0 to 2);
      C440TRCCYCLE         : out std_ulogic;
      C440TRCEXECUTIONSTATUS : out std_logic_vector(0 to 4);
      C440TRCTRACESTATUS   : out std_logic_vector(0 to 6);
      C440TRCTRIGGEREVENTOUT : out std_ulogic;
      C440TRCTRIGGEREVENTTYPE : out std_logic_vector(0 to 13);
      DMA0LLRSTENGINEACK   : out std_ulogic;
      DMA0LLRXDSTRDYN      : out std_ulogic;
      DMA0LLTXD            : out std_logic_vector(0 to 31);
      DMA0LLTXEOFN         : out std_ulogic;
      DMA0LLTXEOPN         : out std_ulogic;
      DMA0LLTXREM          : out std_logic_vector(0 to 3);
      DMA0LLTXSOFN         : out std_ulogic;
      DMA0LLTXSOPN         : out std_ulogic;
      DMA0LLTXSRCRDYN      : out std_ulogic;
      DMA0RXIRQ            : out std_ulogic;
      DMA0TXIRQ            : out std_ulogic;
      DMA1LLRSTENGINEACK   : out std_ulogic;
      DMA1LLRXDSTRDYN      : out std_ulogic;
      DMA1LLTXD            : out std_logic_vector(0 to 31);
      DMA1LLTXEOFN         : out std_ulogic;
      DMA1LLTXEOPN         : out std_ulogic;
      DMA1LLTXREM          : out std_logic_vector(0 to 3);
      DMA1LLTXSOFN         : out std_ulogic;
      DMA1LLTXSOPN         : out std_ulogic;
      DMA1LLTXSRCRDYN      : out std_ulogic;
      DMA1RXIRQ            : out std_ulogic;
      DMA1TXIRQ            : out std_ulogic;
      DMA2LLRSTENGINEACK   : out std_ulogic;
      DMA2LLRXDSTRDYN      : out std_ulogic;
      DMA2LLTXD            : out std_logic_vector(0 to 31);
      DMA2LLTXEOFN         : out std_ulogic;
      DMA2LLTXEOPN         : out std_ulogic;
      DMA2LLTXREM          : out std_logic_vector(0 to 3);
      DMA2LLTXSOFN         : out std_ulogic;
      DMA2LLTXSOPN         : out std_ulogic;
      DMA2LLTXSRCRDYN      : out std_ulogic;
      DMA2RXIRQ            : out std_ulogic;
      DMA2TXIRQ            : out std_ulogic;
      DMA3LLRSTENGINEACK   : out std_ulogic;
      DMA3LLRXDSTRDYN      : out std_ulogic;
      DMA3LLTXD            : out std_logic_vector(0 to 31);
      DMA3LLTXEOFN         : out std_ulogic;
      DMA3LLTXEOPN         : out std_ulogic;
      DMA3LLTXREM          : out std_logic_vector(0 to 3);
      DMA3LLTXSOFN         : out std_ulogic;
      DMA3LLTXSOPN         : out std_ulogic;
      DMA3LLTXSRCRDYN      : out std_ulogic;
      DMA3RXIRQ            : out std_ulogic;
      DMA3TXIRQ            : out std_ulogic;
      MIMCADDRESS          : out std_logic_vector(0 to 35);
      MIMCADDRESSVALID     : out std_ulogic;
      MIMCBANKCONFLICT     : out std_ulogic;
      MIMCBYTEENABLE       : out std_logic_vector(0 to 15);
      MIMCREADNOTWRITE     : out std_ulogic;
      MIMCROWCONFLICT      : out std_ulogic;
      MIMCWRITEDATA        : out std_logic_vector(0 to 127);
      MIMCWRITEDATAVALID   : out std_ulogic;
      PPCCPMINTERCONNECTBUSY : out std_ulogic;
      PPCDMDCRABUS         : out std_logic_vector(0 to 9);
      PPCDMDCRDBUSOUT      : out std_logic_vector(0 to 31);
      PPCDMDCRREAD         : out std_ulogic;
      PPCDMDCRUABUS        : out std_logic_vector(20 to 21);
      PPCDMDCRWRITE        : out std_ulogic;
      PPCDSDCRACK          : out std_ulogic;
      PPCDSDCRDBUSIN       : out std_logic_vector(0 to 31);
      PPCDSDCRTIMEOUTWAIT  : out std_ulogic;
      PPCEICINTERCONNECTIRQ : out std_ulogic;
      PPCMPLBABORT         : out std_ulogic;
      PPCMPLBABUS          : out std_logic_vector(0 to 31);
      PPCMPLBBE            : out std_logic_vector(0 to 15);
      PPCMPLBBUSLOCK       : out std_ulogic;
      PPCMPLBLOCKERR       : out std_ulogic;
      PPCMPLBPRIORITY      : out std_logic_vector(0 to 1);
      PPCMPLBRDBURST       : out std_ulogic;
      PPCMPLBREQUEST       : out std_ulogic;
      PPCMPLBRNW           : out std_ulogic;
      PPCMPLBSIZE          : out std_logic_vector(0 to 3);
      PPCMPLBTATTRIBUTE    : out std_logic_vector(0 to 15);
      PPCMPLBTYPE          : out std_logic_vector(0 to 2);
      PPCMPLBUABUS         : out std_logic_vector(28 to 31);
      PPCMPLBWRBURST       : out std_ulogic;
      PPCMPLBWRDBUS        : out std_logic_vector(0 to 127);
      PPCS0PLBADDRACK      : out std_ulogic;
      PPCS0PLBMBUSY        : out std_logic_vector(0 to 3);
      PPCS0PLBMIRQ         : out std_logic_vector(0 to 3);
      PPCS0PLBMRDERR       : out std_logic_vector(0 to 3);
      PPCS0PLBMWRERR       : out std_logic_vector(0 to 3);
      PPCS0PLBRDBTERM      : out std_ulogic;
      PPCS0PLBRDCOMP       : out std_ulogic;
      PPCS0PLBRDDACK       : out std_ulogic;
      PPCS0PLBRDDBUS       : out std_logic_vector(0 to 127);
      PPCS0PLBRDWDADDR     : out std_logic_vector(0 to 3);
      PPCS0PLBREARBITRATE  : out std_ulogic;
      PPCS0PLBSSIZE        : out std_logic_vector(0 to 1);
      PPCS0PLBWAIT         : out std_ulogic;
      PPCS0PLBWRBTERM      : out std_ulogic;
      PPCS0PLBWRCOMP       : out std_ulogic;
      PPCS0PLBWRDACK       : out std_ulogic;
      PPCS1PLBADDRACK      : out std_ulogic;
      PPCS1PLBMBUSY        : out std_logic_vector(0 to 3);
      PPCS1PLBMIRQ         : out std_logic_vector(0 to 3);
      PPCS1PLBMRDERR       : out std_logic_vector(0 to 3);
      PPCS1PLBMWRERR       : out std_logic_vector(0 to 3);
      PPCS1PLBRDBTERM      : out std_ulogic;
      PPCS1PLBRDCOMP       : out std_ulogic;
      PPCS1PLBRDDACK       : out std_ulogic;
      PPCS1PLBRDDBUS       : out std_logic_vector(0 to 127);
      PPCS1PLBRDWDADDR     : out std_logic_vector(0 to 3);
      PPCS1PLBREARBITRATE  : out std_ulogic;
      PPCS1PLBSSIZE        : out std_logic_vector(0 to 1);
      PPCS1PLBWAIT         : out std_ulogic;
      PPCS1PLBWRBTERM      : out std_ulogic;
      PPCS1PLBWRCOMP       : out std_ulogic;
      PPCS1PLBWRDACK       : out std_ulogic;

      CPMC440CLK           : in std_ulogic;
      CPMC440CLKEN         : in std_ulogic;
      CPMC440CORECLOCKINACTIVE : in std_ulogic;
      CPMC440TIMERCLOCK    : in std_ulogic;
      CPMDCRCLK            : in std_ulogic;
      CPMDMA0LLCLK         : in std_ulogic;
      CPMDMA1LLCLK         : in std_ulogic;
      CPMDMA2LLCLK         : in std_ulogic;
      CPMDMA3LLCLK         : in std_ulogic;
      CPMFCMCLK            : in std_ulogic;
      CPMINTERCONNECTCLK   : in std_ulogic;
      CPMINTERCONNECTCLKEN : in std_ulogic;
      CPMINTERCONNECTCLKNTO1 : in std_ulogic;
      CPMMCCLK             : in std_ulogic;
      CPMPPCMPLBCLK        : in std_ulogic;
      CPMPPCS0PLBCLK       : in std_ulogic;
      CPMPPCS1PLBCLK       : in std_ulogic;
      DBGC440DEBUGHALT     : in std_ulogic;
      DBGC440SYSTEMSTATUS  : in std_logic_vector(0 to 4);
      DBGC440UNCONDDEBUGEVENT : in std_ulogic;
      DCRPPCDMACK          : in std_ulogic;
      DCRPPCDMDBUSIN       : in std_logic_vector(0 to 31);
      DCRPPCDMTIMEOUTWAIT  : in std_ulogic;
      DCRPPCDSABUS         : in std_logic_vector(0 to 9);
      DCRPPCDSDBUSOUT      : in std_logic_vector(0 to 31);
      DCRPPCDSREAD         : in std_ulogic;
      DCRPPCDSWRITE        : in std_ulogic;
      EICC440CRITIRQ       : in std_ulogic;
      EICC440EXTIRQ        : in std_ulogic;
      FCMAPUCONFIRMINSTR   : in std_ulogic;
      FCMAPUCR             : in std_logic_vector(0 to 3);
      FCMAPUDONE           : in std_ulogic;
      FCMAPUEXCEPTION      : in std_ulogic;
      FCMAPUFPSCRFEX       : in std_ulogic;
      FCMAPURESULT         : in std_logic_vector(0 to 31);
      FCMAPURESULTVALID    : in std_ulogic;
      FCMAPUSLEEPNOTREADY  : in std_ulogic;
      FCMAPUSTOREDATA      : in std_logic_vector(0 to 127);
      GSR                  : in std_ulogic;
      JTGC440TCK           : in std_ulogic;
      JTGC440TDI           : in std_ulogic;
      JTGC440TMS           : in std_ulogic;
      JTGC440TRSTNEG       : in std_ulogic;
      LLDMA0RSTENGINEREQ   : in std_ulogic;
      LLDMA0RXD            : in std_logic_vector(0 to 31);
      LLDMA0RXEOFN         : in std_ulogic;
      LLDMA0RXEOPN         : in std_ulogic;
      LLDMA0RXREM          : in std_logic_vector(0 to 3);
      LLDMA0RXSOFN         : in std_ulogic;
      LLDMA0RXSOPN         : in std_ulogic;
      LLDMA0RXSRCRDYN      : in std_ulogic;
      LLDMA0TXDSTRDYN      : in std_ulogic;
      LLDMA1RSTENGINEREQ   : in std_ulogic;
      LLDMA1RXD            : in std_logic_vector(0 to 31);
      LLDMA1RXEOFN         : in std_ulogic;
      LLDMA1RXEOPN         : in std_ulogic;
      LLDMA1RXREM          : in std_logic_vector(0 to 3);
      LLDMA1RXSOFN         : in std_ulogic;
      LLDMA1RXSOPN         : in std_ulogic;
      LLDMA1RXSRCRDYN      : in std_ulogic;
      LLDMA1TXDSTRDYN      : in std_ulogic;
      LLDMA2RSTENGINEREQ   : in std_ulogic;
      LLDMA2RXD            : in std_logic_vector(0 to 31);
      LLDMA2RXEOFN         : in std_ulogic;
      LLDMA2RXEOPN         : in std_ulogic;
      LLDMA2RXREM          : in std_logic_vector(0 to 3);
      LLDMA2RXSOFN         : in std_ulogic;
      LLDMA2RXSOPN         : in std_ulogic;
      LLDMA2RXSRCRDYN      : in std_ulogic;
      LLDMA2TXDSTRDYN      : in std_ulogic;
      LLDMA3RSTENGINEREQ   : in std_ulogic;
      LLDMA3RXD            : in std_logic_vector(0 to 31);
      LLDMA3RXEOFN         : in std_ulogic;
      LLDMA3RXEOPN         : in std_ulogic;
      LLDMA3RXREM          : in std_logic_vector(0 to 3);
      LLDMA3RXSOFN         : in std_ulogic;
      LLDMA3RXSOPN         : in std_ulogic;
      LLDMA3RXSRCRDYN      : in std_ulogic;
      LLDMA3TXDSTRDYN      : in std_ulogic;
      MCMIADDRREADYTOACCEPT : in std_ulogic;
      MCMIREADDATA         : in std_logic_vector(0 to 127);
      MCMIREADDATAERR      : in std_ulogic;
      MCMIREADDATAVALID    : in std_ulogic;
      PLBPPCMADDRACK       : in std_ulogic;
      PLBPPCMMBUSY         : in std_ulogic;
      PLBPPCMMIRQ          : in std_ulogic;
      PLBPPCMMRDERR        : in std_ulogic;
      PLBPPCMMWRERR        : in std_ulogic;
      PLBPPCMRDBTERM       : in std_ulogic;
      PLBPPCMRDDACK        : in std_ulogic;
      PLBPPCMRDDBUS        : in std_logic_vector(0 to 127);
      PLBPPCMRDPENDPRI     : in std_logic_vector(0 to 1);
      PLBPPCMRDPENDREQ     : in std_ulogic;
      PLBPPCMRDWDADDR      : in std_logic_vector(0 to 3);
      PLBPPCMREARBITRATE   : in std_ulogic;
      PLBPPCMREQPRI        : in std_logic_vector(0 to 1);
      PLBPPCMSSIZE         : in std_logic_vector(0 to 1);
      PLBPPCMTIMEOUT       : in std_ulogic;
      PLBPPCMWRBTERM       : in std_ulogic;
      PLBPPCMWRDACK        : in std_ulogic;
      PLBPPCMWRPENDPRI     : in std_logic_vector(0 to 1);
      PLBPPCMWRPENDREQ     : in std_ulogic;
      PLBPPCS0ABORT        : in std_ulogic;
      PLBPPCS0ABUS         : in std_logic_vector(0 to 31);
      PLBPPCS0BE           : in std_logic_vector(0 to 15);
      PLBPPCS0BUSLOCK      : in std_ulogic;
      PLBPPCS0LOCKERR      : in std_ulogic;
      PLBPPCS0MASTERID     : in std_logic_vector(0 to 1);
      PLBPPCS0MSIZE        : in std_logic_vector(0 to 1);
      PLBPPCS0PAVALID      : in std_ulogic;
      PLBPPCS0RDBURST      : in std_ulogic;
      PLBPPCS0RDPENDPRI    : in std_logic_vector(0 to 1);
      PLBPPCS0RDPENDREQ    : in std_ulogic;
      PLBPPCS0RDPRIM       : in std_ulogic;
      PLBPPCS0REQPRI       : in std_logic_vector(0 to 1);
      PLBPPCS0RNW          : in std_ulogic;
      PLBPPCS0SAVALID      : in std_ulogic;
      PLBPPCS0SIZE         : in std_logic_vector(0 to 3);
      PLBPPCS0TATTRIBUTE   : in std_logic_vector(0 to 15);
      PLBPPCS0TYPE         : in std_logic_vector(0 to 2);
      PLBPPCS0UABUS        : in std_logic_vector(28 to 31);
      PLBPPCS0WRBURST      : in std_ulogic;
      PLBPPCS0WRDBUS       : in std_logic_vector(0 to 127);
      PLBPPCS0WRPENDPRI    : in std_logic_vector(0 to 1);
      PLBPPCS0WRPENDREQ    : in std_ulogic;
      PLBPPCS0WRPRIM       : in std_ulogic;
      PLBPPCS1ABORT        : in std_ulogic;
      PLBPPCS1ABUS         : in std_logic_vector(0 to 31);
      PLBPPCS1BE           : in std_logic_vector(0 to 15);
      PLBPPCS1BUSLOCK      : in std_ulogic;
      PLBPPCS1LOCKERR      : in std_ulogic;
      PLBPPCS1MASTERID     : in std_logic_vector(0 to 1);
      PLBPPCS1MSIZE        : in std_logic_vector(0 to 1);
      PLBPPCS1PAVALID      : in std_ulogic;
      PLBPPCS1RDBURST      : in std_ulogic;
      PLBPPCS1RDPENDPRI    : in std_logic_vector(0 to 1);
      PLBPPCS1RDPENDREQ    : in std_ulogic;
      PLBPPCS1RDPRIM       : in std_ulogic;
      PLBPPCS1REQPRI       : in std_logic_vector(0 to 1);
      PLBPPCS1RNW          : in std_ulogic;
      PLBPPCS1SAVALID      : in std_ulogic;
      PLBPPCS1SIZE         : in std_logic_vector(0 to 3);
      PLBPPCS1TATTRIBUTE   : in std_logic_vector(0 to 15);
      PLBPPCS1TYPE         : in std_logic_vector(0 to 2);
      PLBPPCS1UABUS        : in std_logic_vector(28 to 31);
      PLBPPCS1WRBURST      : in std_ulogic;
      PLBPPCS1WRDBUS       : in std_logic_vector(0 to 127);
      PLBPPCS1WRPENDPRI    : in std_logic_vector(0 to 1);
      PLBPPCS1WRPENDREQ    : in std_ulogic;
      PLBPPCS1WRPRIM       : in std_ulogic;
      RSTC440RESETCHIP     : in std_ulogic;
      RSTC440RESETCORE     : in std_ulogic;
      RSTC440RESETSYSTEM   : in std_ulogic;
      TIEC440DCURDLDCACHEPLBPRIO : in std_logic_vector(0 to 1);
      TIEC440DCURDNONCACHEPLBPRIO : in std_logic_vector(0 to 1);
      TIEC440DCURDTOUCHPLBPRIO : in std_logic_vector(0 to 1);
      TIEC440DCURDURGENTPLBPRIO : in std_logic_vector(0 to 1);
      TIEC440DCUWRFLUSHPLBPRIO : in std_logic_vector(0 to 1);
      TIEC440DCUWRSTOREPLBPRIO : in std_logic_vector(0 to 1);
      TIEC440DCUWRURGENTPLBPRIO : in std_logic_vector(0 to 1);
      TIEC440ENDIANRESET   : in std_ulogic;
      TIEC440ERPNRESET     : in std_logic_vector(0 to 3);
      TIEC440ICURDFETCHPLBPRIO : in std_logic_vector(0 to 1);
      TIEC440ICURDSPECPLBPRIO : in std_logic_vector(0 to 1);
      TIEC440ICURDTOUCHPLBPRIO : in std_logic_vector(0 to 1);
      TIEC440PIR           : in std_logic_vector(28 to 31);
      TIEC440PVR           : in std_logic_vector(28 to 31);
      TIEC440USERRESET     : in std_logic_vector(0 to 3);
      TIEDCRBASEADDR       : in std_logic_vector(0 to 1);
      TRCC440TRACEDISABLE  : in std_ulogic;
      TRCC440TRIGGEREVENTIN : in std_ulogic;

      APU_CONTROL          : in std_logic_vector(0 to 16);
      APU_UDI0             : in std_logic_vector(0 to 23);
      APU_UDI1             : in std_logic_vector(0 to 23);
      APU_UDI10            : in std_logic_vector(0 to 23);
      APU_UDI11            : in std_logic_vector(0 to 23);
      APU_UDI12            : in std_logic_vector(0 to 23);
      APU_UDI13            : in std_logic_vector(0 to 23);
      APU_UDI14            : in std_logic_vector(0 to 23);
      APU_UDI15            : in std_logic_vector(0 to 23);
      APU_UDI2             : in std_logic_vector(0 to 23);
      APU_UDI3             : in std_logic_vector(0 to 23);
      APU_UDI4             : in std_logic_vector(0 to 23);
      APU_UDI5             : in std_logic_vector(0 to 23);
      APU_UDI6             : in std_logic_vector(0 to 23);
      APU_UDI7             : in std_logic_vector(0 to 23);
      APU_UDI8             : in std_logic_vector(0 to 23);
      APU_UDI9             : in std_logic_vector(0 to 23);
--      CLOCK_DELAY          : in std_ulogic;
      CLOCK_DELAY          : in std_logic_vector(0 to 4);
      DCR_AUTOLOCK_ENABLE  : in std_ulogic;
      DMA0_CONTROL         : in std_logic_vector(0 to 7);
      DMA0_RXCHANNELCTRL   : in std_logic_vector(0 to 31);
      DMA0_RXIRQTIMER      : in std_logic_vector(0 to 9);
      DMA0_TXCHANNELCTRL   : in std_logic_vector(0 to 31);
      DMA0_TXIRQTIMER      : in std_logic_vector(0 to 9);
      DMA1_CONTROL         : in std_logic_vector(0 to 7);
      DMA1_RXCHANNELCTRL   : in std_logic_vector(0 to 31);
      DMA1_RXIRQTIMER      : in std_logic_vector(0 to 9);
      DMA1_TXCHANNELCTRL   : in std_logic_vector(0 to 31);
      DMA1_TXIRQTIMER      : in std_logic_vector(0 to 9);
      DMA2_CONTROL         : in std_logic_vector(0 to 7);
      DMA2_RXCHANNELCTRL   : in std_logic_vector(0 to 31);
      DMA2_RXIRQTIMER      : in std_logic_vector(0 to 9);
      DMA2_TXCHANNELCTRL   : in std_logic_vector(0 to 31);
      DMA2_TXIRQTIMER      : in std_logic_vector(0 to 9);
      DMA3_CONTROL         : in std_logic_vector(0 to 7);
      DMA3_RXCHANNELCTRL   : in std_logic_vector(0 to 31);
      DMA3_RXIRQTIMER      : in std_logic_vector(0 to 9);
      DMA3_TXCHANNELCTRL   : in std_logic_vector(0 to 31);
      DMA3_TXIRQTIMER      : in std_logic_vector(0 to 9);
      INTERCONNECT_IMASK   : in std_logic_vector(0 to 31);
      INTERCONNECT_TMPL_SEL : in std_logic_vector(0 to 31);
      MI_ARBCONFIG         : in std_logic_vector(0 to 31);
      MI_BANKCONFLICT_MASK : in std_logic_vector(0 to 31);
      MI_CONTROL           : in std_logic_vector(0 to 31);
      MI_ROWCONFLICT_MASK  : in std_logic_vector(0 to 31);
      PPCDM_ASYNCMODE      : in std_ulogic;
      PPCDS_ASYNCMODE      : in std_ulogic;
      PPCM_ARBCONFIG       : in std_logic_vector(0 to 31);
      PPCM_CONTROL         : in std_logic_vector(0 to 31);
      PPCM_COUNTER         : in std_logic_vector(0 to 31);
      PPCS0_ADDRMAP_TMPL0  : in std_logic_vector(0 to 31);
      PPCS0_ADDRMAP_TMPL1  : in std_logic_vector(0 to 31);
      PPCS0_ADDRMAP_TMPL2  : in std_logic_vector(0 to 31);
      PPCS0_ADDRMAP_TMPL3  : in std_logic_vector(0 to 31);
      PPCS0_CONTROL        : in std_logic_vector(0 to 31);
      PPCS0_WIDTH_128N64   : in std_ulogic;
      PPCS1_ADDRMAP_TMPL0  : in std_logic_vector(0 to 31);
      PPCS1_ADDRMAP_TMPL1  : in std_logic_vector(0 to 31);
      PPCS1_ADDRMAP_TMPL2  : in std_logic_vector(0 to 31);
      PPCS1_ADDRMAP_TMPL3  : in std_logic_vector(0 to 31);
      PPCS1_CONTROL        : in std_logic_vector(0 to 31);
      PPCS1_WIDTH_128N64   : in std_ulogic;
      XBAR_ADDRMAP_TMPL0   : in std_logic_vector(0 to 31);
      XBAR_ADDRMAP_TMPL1   : in std_logic_vector(0 to 31);
      XBAR_ADDRMAP_TMPL2   : in std_logic_vector(0 to 31);
      XBAR_ADDRMAP_TMPL3   : in std_logic_vector(0 to 31)
    );
  end component;

	constant IN_DELAY : time :=  1 ps;
	constant OUT_DELAY : time := 0 ps;
	constant CLK_DELAY : time := 0 ps;
  	constant ZERO_DELAY : time := 0 ps;

	constant PATH_DELAY : VitalDelayType01 := (100 ps, 100 ps);


	signal   DMA3_TXCHANNELCTRL_BINARY  :  std_logic_vector(0 to 31) := To_StdLogicVector(DMA3_TXCHANNELCTRL);
	signal   DMA3_CONTROL_BINARY  :  std_logic_vector(0 to 7) := To_StdLogicVector(DMA3_CONTROL);
	signal   DMA3_RXCHANNELCTRL_BINARY  :  std_logic_vector(0 to 31) := To_StdLogicVector(DMA3_RXCHANNELCTRL);
	signal   DMA3_TXIRQTIMER_BINARY  :  std_logic_vector(0 to 9) := To_StdLogicVector(DMA3_TXIRQTIMER)(9 downto 0);
	signal   DMA3_RXIRQTIMER_BINARY  :  std_logic_vector(0 to 9) := To_StdLogicVector(DMA3_RXIRQTIMER)(9 downto 0);
	signal   DMA2_TXCHANNELCTRL_BINARY  :  std_logic_vector(0 to 31) := To_StdLogicVector(DMA2_TXCHANNELCTRL);
	signal   DMA2_CONTROL_BINARY  :  std_logic_vector(0 to 7) := To_StdLogicVector(DMA2_CONTROL);
	signal   DMA2_RXCHANNELCTRL_BINARY  :  std_logic_vector(0 to 31) := To_StdLogicVector(DMA2_RXCHANNELCTRL);
	signal   DMA2_TXIRQTIMER_BINARY  :  std_logic_vector(0 to 9) := To_StdLogicVector(DMA2_TXIRQTIMER)(9 downto 0);
	signal   DMA2_RXIRQTIMER_BINARY  :  std_logic_vector(0 to 9) := To_StdLogicVector(DMA2_RXIRQTIMER)(9 downto 0);
	signal   PPCM_CONTROL_BINARY  :  std_logic_vector(0 to 31) := To_StdLogicVector(PPCM_CONTROL);
	signal   PPCM_COUNTER_BINARY  :  std_logic_vector(0 to 31) := To_StdLogicVector(PPCM_COUNTER);
	signal   PPCM_ARBCONFIG_BINARY  :  std_logic_vector(0 to 31) := To_StdLogicVector(PPCM_ARBCONFIG);
	signal   DMA1_RXIRQTIMER_BINARY  :  std_logic_vector(0 to 9) := To_StdLogicVector(DMA1_RXIRQTIMER)(9 downto 0);
	signal   DMA1_TXIRQTIMER_BINARY  :  std_logic_vector(0 to 9) := To_StdLogicVector(DMA1_TXIRQTIMER)(9 downto 0);
	signal   DMA1_RXCHANNELCTRL_BINARY  :  std_logic_vector(0 to 31) := To_StdLogicVector(DMA1_RXCHANNELCTRL);
	signal   DMA1_CONTROL_BINARY  :  std_logic_vector(0 to 7) := To_StdLogicVector(DMA1_CONTROL);
	signal   DMA1_TXCHANNELCTRL_BINARY  :  std_logic_vector(0 to 31) := To_StdLogicVector(DMA1_TXCHANNELCTRL);
	signal   DMA0_RXIRQTIMER_BINARY  :  std_logic_vector(0 to 9) := To_StdLogicVector(DMA0_RXIRQTIMER)(9 downto 0);
	signal   DMA0_TXIRQTIMER_BINARY  :  std_logic_vector(0 to 9) := To_StdLogicVector(DMA0_TXIRQTIMER)(9 downto 0);
	signal   DMA0_RXCHANNELCTRL_BINARY  :  std_logic_vector(0 to 31) := To_StdLogicVector(DMA0_RXCHANNELCTRL);
	signal   DMA0_CONTROL_BINARY  :  std_logic_vector(0 to 7) := To_StdLogicVector(DMA0_CONTROL);
	signal   DMA0_TXCHANNELCTRL_BINARY  :  std_logic_vector(0 to 31) := To_StdLogicVector(DMA0_TXCHANNELCTRL);
	signal   MI_ROWCONFLICT_MASK_BINARY  :  std_logic_vector(0 to 31) := To_StdLogicVector(MI_ROWCONFLICT_MASK);
	signal   MI_BANKCONFLICT_MASK_BINARY  :  std_logic_vector(0 to 31) := To_StdLogicVector(MI_BANKCONFLICT_MASK);
	signal   MI_ARBCONFIG_BINARY  :  std_logic_vector(0 to 31) := To_StdLogicVector(MI_ARBCONFIG);
	signal   MI_CONTROL_BINARY  :  std_logic_vector(0 to 31) := To_StdLogicVector(MI_CONTROL);
	signal   APU_UDI0_BINARY  :  std_logic_vector(0 to 23) := To_StdLogicVector(APU_UDI0);
	signal   APU_UDI1_BINARY  :  std_logic_vector(0 to 23) := To_StdLogicVector(APU_UDI1);
	signal   APU_UDI2_BINARY  :  std_logic_vector(0 to 23) := To_StdLogicVector(APU_UDI2);
	signal   APU_UDI3_BINARY  :  std_logic_vector(0 to 23) := To_StdLogicVector(APU_UDI3);
	signal   APU_UDI4_BINARY  :  std_logic_vector(0 to 23) := To_StdLogicVector(APU_UDI4);
	signal   APU_UDI5_BINARY  :  std_logic_vector(0 to 23) := To_StdLogicVector(APU_UDI5);
	signal   APU_UDI6_BINARY  :  std_logic_vector(0 to 23) := To_StdLogicVector(APU_UDI6);
	signal   APU_UDI7_BINARY  :  std_logic_vector(0 to 23) := To_StdLogicVector(APU_UDI7);
	signal   APU_UDI8_BINARY  :  std_logic_vector(0 to 23) := To_StdLogicVector(APU_UDI8);
	signal   APU_UDI9_BINARY  :  std_logic_vector(0 to 23) := To_StdLogicVector(APU_UDI9);
	signal   APU_UDI10_BINARY  :  std_logic_vector(0 to 23) := To_StdLogicVector(APU_UDI10);
	signal   APU_UDI11_BINARY  :  std_logic_vector(0 to 23) := To_StdLogicVector(APU_UDI11);
	signal   APU_UDI12_BINARY  :  std_logic_vector(0 to 23) := To_StdLogicVector(APU_UDI12);
	signal   APU_UDI13_BINARY  :  std_logic_vector(0 to 23) := To_StdLogicVector(APU_UDI13);
	signal   APU_UDI14_BINARY  :  std_logic_vector(0 to 23) := To_StdLogicVector(APU_UDI14);
	signal   APU_UDI15_BINARY  :  std_logic_vector(0 to 23) := To_StdLogicVector(APU_UDI15);
	signal   APU_CONTROL_BINARY  :  std_logic_vector(0 to 16) := To_StdLogicVector(APU_CONTROL)(16 downto 0);
	signal   INTERCONNECT_IMASK_BINARY  :  std_logic_vector(0 to 31) := To_StdLogicVector(INTERCONNECT_IMASK);
	signal   XBAR_ADDRMAP_TMPL0_BINARY  :  std_logic_vector(0 to 31) := To_StdLogicVector(XBAR_ADDRMAP_TMPL0);
	signal   XBAR_ADDRMAP_TMPL1_BINARY  :  std_logic_vector(0 to 31) := To_StdLogicVector(XBAR_ADDRMAP_TMPL1);
	signal   XBAR_ADDRMAP_TMPL2_BINARY  :  std_logic_vector(0 to 31) := To_StdLogicVector(XBAR_ADDRMAP_TMPL2);
	signal   XBAR_ADDRMAP_TMPL3_BINARY  :  std_logic_vector(0 to 31) := To_StdLogicVector(XBAR_ADDRMAP_TMPL3);
	signal   INTERCONNECT_TMPL_SEL_BINARY  :  std_logic_vector(0 to 31) := To_StdLogicVector(INTERCONNECT_TMPL_SEL);
	signal   PPCS0_CONTROL_BINARY  :  std_logic_vector(0 to 31) := To_StdLogicVector(PPCS0_CONTROL);
	signal   PPCS0_WIDTH_128N64_BINARY  :  std_ulogic;
	signal   PPCS0_ADDRMAP_TMPL0_BINARY  :  std_logic_vector(0 to 31) := To_StdLogicVector(PPCS0_ADDRMAP_TMPL0);
	signal   PPCS0_ADDRMAP_TMPL1_BINARY  :  std_logic_vector(0 to 31) := To_StdLogicVector(PPCS0_ADDRMAP_TMPL1);
	signal   PPCS0_ADDRMAP_TMPL2_BINARY  :  std_logic_vector(0 to 31) := To_StdLogicVector(PPCS0_ADDRMAP_TMPL2);
	signal   PPCS0_ADDRMAP_TMPL3_BINARY  :  std_logic_vector(0 to 31) := To_StdLogicVector(PPCS0_ADDRMAP_TMPL3);
	signal   PPCS1_CONTROL_BINARY  :  std_logic_vector(0 to 31) := To_StdLogicVector(PPCS1_CONTROL);
	signal   PPCS1_WIDTH_128N64_BINARY  :  std_ulogic;
	signal   PPCS1_ADDRMAP_TMPL0_BINARY  :  std_logic_vector(0 to 31) := To_StdLogicVector(PPCS1_ADDRMAP_TMPL0);
	signal   PPCS1_ADDRMAP_TMPL1_BINARY  :  std_logic_vector(0 to 31) := To_StdLogicVector(PPCS1_ADDRMAP_TMPL1);
	signal   PPCS1_ADDRMAP_TMPL2_BINARY  :  std_logic_vector(0 to 31) := To_StdLogicVector(PPCS1_ADDRMAP_TMPL2);
	signal   PPCS1_ADDRMAP_TMPL3_BINARY  :  std_logic_vector(0 to 31) := To_StdLogicVector(PPCS1_ADDRMAP_TMPL3);
	signal   PPCDM_ASYNCMODE_BINARY  :  std_ulogic;
	signal   PPCDS_ASYNCMODE_BINARY  :  std_ulogic;
	signal   DCR_AUTOLOCK_ENABLE_BINARY  :  std_ulogic;
	signal   CLOCK_DELAY_BINARY  :   std_logic_vector(0 to 4);

	signal   DMA0LLRSTENGINEACK_out  :  std_ulogic;
	signal   DMA0LLRXDSTRDYN_out  :  std_ulogic;
	signal   DMA0LLTXD_out  :  std_logic_vector(0 to 31);
	signal   DMA0LLTXEOFN_out  :  std_ulogic;
	signal   DMA0LLTXEOPN_out  :  std_ulogic;
	signal   DMA0LLTXREM_out  :  std_logic_vector(0 to 3);
	signal   DMA0LLTXSOFN_out  :  std_ulogic;
	signal   DMA0LLTXSOPN_out  :  std_ulogic;
	signal   DMA0LLTXSRCRDYN_out  :  std_ulogic;
	signal   DMA0RXIRQ_out  :  std_ulogic;
	signal   DMA0TXIRQ_out  :  std_ulogic;
	signal   DMA1LLRSTENGINEACK_out  :  std_ulogic;
	signal   DMA1LLRXDSTRDYN_out  :  std_ulogic;
	signal   DMA1LLTXD_out  :  std_logic_vector(0 to 31);
	signal   DMA1LLTXEOFN_out  :  std_ulogic;
	signal   DMA1LLTXEOPN_out  :  std_ulogic;
	signal   DMA1LLTXREM_out  :  std_logic_vector(0 to 3);
	signal   DMA1LLTXSOFN_out  :  std_ulogic;
	signal   DMA1LLTXSOPN_out  :  std_ulogic;
	signal   DMA1LLTXSRCRDYN_out  :  std_ulogic;
	signal   DMA1RXIRQ_out  :  std_ulogic;
	signal   DMA1TXIRQ_out  :  std_ulogic;
	signal   DMA2LLRSTENGINEACK_out  :  std_ulogic;
	signal   DMA2LLRXDSTRDYN_out  :  std_ulogic;
	signal   DMA2LLTXD_out  :  std_logic_vector(0 to 31);
	signal   DMA2LLTXEOFN_out  :  std_ulogic;
	signal   DMA2LLTXEOPN_out  :  std_ulogic;
	signal   DMA2LLTXREM_out  :  std_logic_vector(0 to 3);
	signal   DMA2LLTXSOFN_out  :  std_ulogic;
	signal   DMA2LLTXSOPN_out  :  std_ulogic;
	signal   DMA2LLTXSRCRDYN_out  :  std_ulogic;
	signal   DMA2RXIRQ_out  :  std_ulogic;
	signal   DMA2TXIRQ_out  :  std_ulogic;
	signal   DMA3LLRSTENGINEACK_out  :  std_ulogic;
	signal   DMA3LLRXDSTRDYN_out  :  std_ulogic;
	signal   DMA3LLTXD_out  :  std_logic_vector(0 to 31);
	signal   DMA3LLTXEOFN_out  :  std_ulogic;
	signal   DMA3LLTXEOPN_out  :  std_ulogic;
	signal   DMA3LLTXREM_out  :  std_logic_vector(0 to 3);
	signal   DMA3LLTXSOFN_out  :  std_ulogic;
	signal   DMA3LLTXSOPN_out  :  std_ulogic;
	signal   DMA3LLTXSRCRDYN_out  :  std_ulogic;
	signal   DMA3RXIRQ_out  :  std_ulogic;
	signal   DMA3TXIRQ_out  :  std_ulogic;
	signal   PPCDMDCRABUS_out  :  std_logic_vector(0 to 9);
	signal   PPCDMDCRDBUSOUT_out  :  std_logic_vector(0 to 31);
	signal   PPCDMDCRREAD_out  :  std_ulogic;
	signal   PPCDMDCRUABUS_out  :  std_logic_vector(20 to 21);
	signal   PPCDMDCRWRITE_out  :  std_ulogic;
	signal   PPCMPLBABORT_out  :  std_ulogic;
	signal   PPCMPLBABUS_out  :  std_logic_vector(0 to 31);
	signal   PPCMPLBBE_out  :  std_logic_vector(0 to 15);
	signal   PPCMPLBBUSLOCK_out  :  std_ulogic;
	signal   PPCMPLBLOCKERR_out  :  std_ulogic;
	signal   PPCMPLBPRIORITY_out  :  std_logic_vector(0 to 1);
	signal   PPCMPLBRDBURST_out  :  std_ulogic;
	signal   PPCMPLBREQUEST_out  :  std_ulogic;
	signal   PPCMPLBRNW_out  :  std_ulogic;
	signal   PPCMPLBSIZE_out  :  std_logic_vector(0 to 3);
	signal   PPCMPLBTATTRIBUTE_out  :  std_logic_vector(0 to 15);
	signal   PPCMPLBTYPE_out  :  std_logic_vector(0 to 2);
	signal   PPCMPLBUABUS_out  :  std_logic_vector(28 to 31);
	signal   PPCMPLBWRBURST_out  :  std_ulogic;
	signal   PPCMPLBWRDBUS_out  :  std_logic_vector(0 to 127);
	signal   PPCS0PLBADDRACK_out  :  std_ulogic;
	signal   PPCS0PLBMBUSY_out  :  std_logic_vector(0 to 3);
	signal   PPCS0PLBMIRQ_out  :  std_logic_vector(0 to 3);
	signal   PPCS0PLBMRDERR_out  :  std_logic_vector(0 to 3);
	signal   PPCS0PLBMWRERR_out  :  std_logic_vector(0 to 3);
	signal   PPCS0PLBRDBTERM_out  :  std_ulogic;
	signal   PPCS0PLBRDCOMP_out  :  std_ulogic;
	signal   PPCS0PLBRDDACK_out  :  std_ulogic;
	signal   PPCS0PLBRDDBUS_out  :  std_logic_vector(0 to 127);
	signal   PPCS0PLBRDWDADDR_out  :  std_logic_vector(0 to 3);
	signal   PPCS0PLBREARBITRATE_out  :  std_ulogic;
	signal   PPCS0PLBSSIZE_out  :  std_logic_vector(0 to 1);
	signal   PPCS0PLBWAIT_out  :  std_ulogic;
	signal   PPCS0PLBWRBTERM_out  :  std_ulogic;
	signal   PPCS0PLBWRCOMP_out  :  std_ulogic;
	signal   PPCS0PLBWRDACK_out  :  std_ulogic;
	signal   PPCS1PLBADDRACK_out  :  std_ulogic;
	signal   PPCS1PLBMBUSY_out  :  std_logic_vector(0 to 3);
	signal   PPCS1PLBMIRQ_out  :  std_logic_vector(0 to 3);
	signal   PPCS1PLBMRDERR_out  :  std_logic_vector(0 to 3);
	signal   PPCS1PLBMWRERR_out  :  std_logic_vector(0 to 3);
	signal   PPCS1PLBRDBTERM_out  :  std_ulogic;
	signal   PPCS1PLBRDCOMP_out  :  std_ulogic;
	signal   PPCS1PLBRDDACK_out  :  std_ulogic;
	signal   PPCS1PLBRDDBUS_out  :  std_logic_vector(0 to 127);
	signal   PPCS1PLBRDWDADDR_out  :  std_logic_vector(0 to 3);
	signal   PPCS1PLBREARBITRATE_out  :  std_ulogic;
	signal   PPCS1PLBSSIZE_out  :  std_logic_vector(0 to 1);
	signal   PPCS1PLBWAIT_out  :  std_ulogic;
	signal   PPCS1PLBWRBTERM_out  :  std_ulogic;
	signal   PPCS1PLBWRCOMP_out  :  std_ulogic;
	signal   PPCS1PLBWRDACK_out  :  std_ulogic;
	signal   APUFCMDECFPUOP_out  :  std_ulogic;
	signal   APUFCMDECLDSTXFERSIZE_out  :  std_logic_vector(0 to 2);
	signal   APUFCMDECLOAD_out  :  std_ulogic;
	signal   APUFCMDECNONAUTON_out  :  std_ulogic;
	signal   APUFCMDECSTORE_out  :  std_ulogic;
	signal   APUFCMDECUDI_out  :  std_logic_vector(0 to 3);
	signal   APUFCMDECUDIVALID_out  :  std_ulogic;
	signal   APUFCMENDIAN_out  :  std_ulogic;
	signal   APUFCMFLUSH_out  :  std_ulogic;
	signal   APUFCMINSTRUCTION_out  :  std_logic_vector(0 to 31);
	signal   APUFCMINSTRVALID_out  :  std_ulogic;
	signal   APUFCMLOADBYTEADDR_out  :  std_logic_vector(0 to 3);
	signal   APUFCMLOADDATA_out  :  std_logic_vector(0 to 127);
	signal   APUFCMLOADDVALID_out  :  std_ulogic;
	signal   APUFCMMSRFE0_out  :  std_ulogic;
	signal   APUFCMMSRFE1_out  :  std_ulogic;
	signal   APUFCMNEXTINSTRREADY_out  :  std_ulogic;
	signal   APUFCMOPERANDVALID_out  :  std_ulogic;
	signal   APUFCMRADATA_out  :  std_logic_vector(0 to 31);
	signal   APUFCMRBDATA_out  :  std_logic_vector(0 to 31);
	signal   APUFCMWRITEBACKOK_out  :  std_ulogic;
	signal   C440CPMCORESLEEPREQ_out  :  std_ulogic;
	signal   C440CPMDECIRPTREQ_out  :  std_ulogic;
	signal   C440CPMFITIRPTREQ_out  :  std_ulogic;
	signal   C440CPMMSRCE_out  :  std_ulogic;
	signal   C440CPMMSREE_out  :  std_ulogic;
	signal   C440CPMTIMERRESETREQ_out  :  std_ulogic;
	signal   C440CPMWDIRPTREQ_out  :  std_ulogic;
	signal   C440DBGSYSTEMCONTROL_out  :  std_logic_vector(0 to 7);
	signal   C440JTGTDO_out  :  std_ulogic;
	signal   C440JTGTDOEN_out  :  std_ulogic;
	signal   C440MACHINECHECK_out  :  std_ulogic;
	signal   C440RSTCHIPRESETREQ_out  :  std_ulogic;
	signal   C440RSTCORERESETREQ_out  :  std_ulogic;
	signal   C440RSTSYSTEMRESETREQ_out  :  std_ulogic;
	signal   C440TRCBRANCHSTATUS_out  :  std_logic_vector(0 to 2);
	signal   C440TRCCYCLE_out  :  std_ulogic;
	signal   C440TRCEXECUTIONSTATUS_out  :  std_logic_vector(0 to 4);
	signal   C440TRCTRACESTATUS_out  :  std_logic_vector(0 to 6);
	signal   C440TRCTRIGGEREVENTOUT_out  :  std_ulogic;
	signal   C440TRCTRIGGEREVENTTYPE_out  :  std_logic_vector(0 to 13);
	signal   MIMCADDRESS_out  :  std_logic_vector(0 to 35);
	signal   MIMCADDRESSVALID_out  :  std_ulogic;
	signal   MIMCBANKCONFLICT_out  :  std_ulogic;
	signal   MIMCBYTEENABLE_out  :  std_logic_vector(0 to 15);
	signal   MIMCREADNOTWRITE_out  :  std_ulogic;
	signal   MIMCROWCONFLICT_out  :  std_ulogic;
	signal   MIMCWRITEDATA_out  :  std_logic_vector(0 to 127);
	signal   MIMCWRITEDATAVALID_out  :  std_ulogic;
	signal   PPCCPMINTERCONNECTBUSY_out  :  std_ulogic;
	signal   PPCDSDCRACK_out  :  std_ulogic;
	signal   PPCDSDCRTIMEOUTWAIT_out  :  std_ulogic;
	signal   PPCDSDCRDBUSIN_out  :  std_logic_vector(0 to 31);
	signal   PPCEICINTERCONNECTIRQ_out  :  std_ulogic;


	signal   DMA0LLRSTENGINEACK_outdelay  :  std_ulogic;
	signal   DMA0LLRXDSTRDYN_outdelay  :  std_ulogic;
	signal   DMA0LLTXD_outdelay  :  std_logic_vector(0 to 31);
	signal   DMA0LLTXEOFN_outdelay  :  std_ulogic;
	signal   DMA0LLTXEOPN_outdelay  :  std_ulogic;
	signal   DMA0LLTXREM_outdelay  :  std_logic_vector(0 to 3);
	signal   DMA0LLTXSOFN_outdelay  :  std_ulogic;
	signal   DMA0LLTXSOPN_outdelay  :  std_ulogic;
	signal   DMA0LLTXSRCRDYN_outdelay  :  std_ulogic;
	signal   DMA0RXIRQ_outdelay  :  std_ulogic;
	signal   DMA0TXIRQ_outdelay  :  std_ulogic;
	signal   DMA1LLRSTENGINEACK_outdelay  :  std_ulogic;
	signal   DMA1LLRXDSTRDYN_outdelay  :  std_ulogic;
	signal   DMA1LLTXD_outdelay  :  std_logic_vector(0 to 31);
	signal   DMA1LLTXEOFN_outdelay  :  std_ulogic;
	signal   DMA1LLTXEOPN_outdelay  :  std_ulogic;
	signal   DMA1LLTXREM_outdelay  :  std_logic_vector(0 to 3);
	signal   DMA1LLTXSOFN_outdelay  :  std_ulogic;
	signal   DMA1LLTXSOPN_outdelay  :  std_ulogic;
	signal   DMA1LLTXSRCRDYN_outdelay  :  std_ulogic;
	signal   DMA1RXIRQ_outdelay  :  std_ulogic;
	signal   DMA1TXIRQ_outdelay  :  std_ulogic;
	signal   DMA2LLRSTENGINEACK_outdelay  :  std_ulogic;
	signal   DMA2LLRXDSTRDYN_outdelay  :  std_ulogic;
	signal   DMA2LLTXD_outdelay  :  std_logic_vector(0 to 31);
	signal   DMA2LLTXEOFN_outdelay  :  std_ulogic;
	signal   DMA2LLTXEOPN_outdelay  :  std_ulogic;
	signal   DMA2LLTXREM_outdelay  :  std_logic_vector(0 to 3);
	signal   DMA2LLTXSOFN_outdelay  :  std_ulogic;
	signal   DMA2LLTXSOPN_outdelay  :  std_ulogic;
	signal   DMA2LLTXSRCRDYN_outdelay  :  std_ulogic;
	signal   DMA2RXIRQ_outdelay  :  std_ulogic;
	signal   DMA2TXIRQ_outdelay  :  std_ulogic;
	signal   DMA3LLRSTENGINEACK_outdelay  :  std_ulogic;
	signal   DMA3LLRXDSTRDYN_outdelay  :  std_ulogic;
	signal   DMA3LLTXD_outdelay  :  std_logic_vector(0 to 31);
	signal   DMA3LLTXEOFN_outdelay  :  std_ulogic;
	signal   DMA3LLTXEOPN_outdelay  :  std_ulogic;
	signal   DMA3LLTXREM_outdelay  :  std_logic_vector(0 to 3);
	signal   DMA3LLTXSOFN_outdelay  :  std_ulogic;
	signal   DMA3LLTXSOPN_outdelay  :  std_ulogic;
	signal   DMA3LLTXSRCRDYN_outdelay  :  std_ulogic;
	signal   DMA3RXIRQ_outdelay  :  std_ulogic;
	signal   DMA3TXIRQ_outdelay  :  std_ulogic;
	signal   PPCDMDCRABUS_outdelay  :  std_logic_vector(0 to 9);
	signal   PPCDMDCRDBUSOUT_outdelay  :  std_logic_vector(0 to 31);
	signal   PPCDMDCRREAD_outdelay  :  std_ulogic;
	signal   PPCDMDCRUABUS_outdelay  :  std_logic_vector(20 to 21);
	signal   PPCDMDCRWRITE_outdelay  :  std_ulogic;
	signal   PPCMPLBABORT_outdelay  :  std_ulogic;
	signal   PPCMPLBABUS_outdelay  :  std_logic_vector(0 to 31);
	signal   PPCMPLBBE_outdelay  :  std_logic_vector(0 to 15);
	signal   PPCMPLBBUSLOCK_outdelay  :  std_ulogic;
	signal   PPCMPLBLOCKERR_outdelay  :  std_ulogic;
	signal   PPCMPLBPRIORITY_outdelay  :  std_logic_vector(0 to 1);
	signal   PPCMPLBRDBURST_outdelay  :  std_ulogic;
	signal   PPCMPLBREQUEST_outdelay  :  std_ulogic;
	signal   PPCMPLBRNW_outdelay  :  std_ulogic;
	signal   PPCMPLBSIZE_outdelay  :  std_logic_vector(0 to 3);
	signal   PPCMPLBTATTRIBUTE_outdelay  :  std_logic_vector(0 to 15);
	signal   PPCMPLBTYPE_outdelay  :  std_logic_vector(0 to 2);
	signal   PPCMPLBUABUS_outdelay  :  std_logic_vector(28 to 31);
	signal   PPCMPLBWRBURST_outdelay  :  std_ulogic;
	signal   PPCMPLBWRDBUS_outdelay  :  std_logic_vector(0 to 127);
	signal   PPCS0PLBADDRACK_outdelay  :  std_ulogic;
	signal   PPCS0PLBMBUSY_outdelay  :  std_logic_vector(0 to 3);
	signal   PPCS0PLBMIRQ_outdelay  :  std_logic_vector(0 to 3);
	signal   PPCS0PLBMRDERR_outdelay  :  std_logic_vector(0 to 3);
	signal   PPCS0PLBMWRERR_outdelay  :  std_logic_vector(0 to 3);
	signal   PPCS0PLBRDBTERM_outdelay  :  std_ulogic;
	signal   PPCS0PLBRDCOMP_outdelay  :  std_ulogic;
	signal   PPCS0PLBRDDACK_outdelay  :  std_ulogic;
	signal   PPCS0PLBRDDBUS_outdelay  :  std_logic_vector(0 to 127);
	signal   PPCS0PLBRDWDADDR_outdelay  :  std_logic_vector(0 to 3);
	signal   PPCS0PLBREARBITRATE_outdelay  :  std_ulogic;
	signal   PPCS0PLBSSIZE_outdelay  :  std_logic_vector(0 to 1);
	signal   PPCS0PLBWAIT_outdelay  :  std_ulogic;
	signal   PPCS0PLBWRBTERM_outdelay  :  std_ulogic;
	signal   PPCS0PLBWRCOMP_outdelay  :  std_ulogic;
	signal   PPCS0PLBWRDACK_outdelay  :  std_ulogic;
	signal   PPCS1PLBADDRACK_outdelay  :  std_ulogic;
	signal   PPCS1PLBMBUSY_outdelay  :  std_logic_vector(0 to 3);
	signal   PPCS1PLBMIRQ_outdelay  :  std_logic_vector(0 to 3);
	signal   PPCS1PLBMRDERR_outdelay  :  std_logic_vector(0 to 3);
	signal   PPCS1PLBMWRERR_outdelay  :  std_logic_vector(0 to 3);
	signal   PPCS1PLBRDBTERM_outdelay  :  std_ulogic;
	signal   PPCS1PLBRDCOMP_outdelay  :  std_ulogic;
	signal   PPCS1PLBRDDACK_outdelay  :  std_ulogic;
	signal   PPCS1PLBRDDBUS_outdelay  :  std_logic_vector(0 to 127);
	signal   PPCS1PLBRDWDADDR_outdelay  :  std_logic_vector(0 to 3);
	signal   PPCS1PLBREARBITRATE_outdelay  :  std_ulogic;
	signal   PPCS1PLBSSIZE_outdelay  :  std_logic_vector(0 to 1);
	signal   PPCS1PLBWAIT_outdelay  :  std_ulogic;
	signal   PPCS1PLBWRBTERM_outdelay  :  std_ulogic;
	signal   PPCS1PLBWRCOMP_outdelay  :  std_ulogic;
	signal   PPCS1PLBWRDACK_outdelay  :  std_ulogic;
	signal   APUFCMDECFPUOP_outdelay  :  std_ulogic;
	signal   APUFCMDECLDSTXFERSIZE_outdelay  :  std_logic_vector(0 to 2);
	signal   APUFCMDECLOAD_outdelay  :  std_ulogic;
	signal   APUFCMDECNONAUTON_outdelay  :  std_ulogic;
	signal   APUFCMDECSTORE_outdelay  :  std_ulogic;
	signal   APUFCMDECUDI_outdelay  :  std_logic_vector(0 to 3);
	signal   APUFCMDECUDIVALID_outdelay  :  std_ulogic;
	signal   APUFCMENDIAN_outdelay  :  std_ulogic;
	signal   APUFCMFLUSH_outdelay  :  std_ulogic;
	signal   APUFCMINSTRUCTION_outdelay  :  std_logic_vector(0 to 31);
	signal   APUFCMINSTRVALID_outdelay  :  std_ulogic;
	signal   APUFCMLOADBYTEADDR_outdelay  :  std_logic_vector(0 to 3);
	signal   APUFCMLOADDATA_outdelay  :  std_logic_vector(0 to 127);
	signal   APUFCMLOADDVALID_outdelay  :  std_ulogic;
	signal   APUFCMMSRFE0_outdelay  :  std_ulogic;
	signal   APUFCMMSRFE1_outdelay  :  std_ulogic;
	signal   APUFCMNEXTINSTRREADY_outdelay  :  std_ulogic;
	signal   APUFCMOPERANDVALID_outdelay  :  std_ulogic;
	signal   APUFCMRADATA_outdelay  :  std_logic_vector(0 to 31);
	signal   APUFCMRBDATA_outdelay  :  std_logic_vector(0 to 31);
	signal   APUFCMWRITEBACKOK_outdelay  :  std_ulogic;
	signal   C440CPMCORESLEEPREQ_outdelay  :  std_ulogic;
	signal   C440CPMDECIRPTREQ_outdelay  :  std_ulogic;
	signal   C440CPMFITIRPTREQ_outdelay  :  std_ulogic;
	signal   C440CPMMSRCE_outdelay  :  std_ulogic;
	signal   C440CPMMSREE_outdelay  :  std_ulogic;
	signal   C440CPMTIMERRESETREQ_outdelay  :  std_ulogic;
	signal   C440CPMWDIRPTREQ_outdelay  :  std_ulogic;
	signal   C440DBGSYSTEMCONTROL_outdelay  :  std_logic_vector(0 to 7);
	signal   C440JTGTDO_outdelay  :  std_ulogic;
	signal   C440JTGTDOEN_outdelay  :  std_ulogic;
	signal   C440MACHINECHECK_outdelay  :  std_ulogic;
	signal   C440RSTCHIPRESETREQ_outdelay  :  std_ulogic;
	signal   C440RSTCORERESETREQ_outdelay  :  std_ulogic;
	signal   C440RSTSYSTEMRESETREQ_outdelay  :  std_ulogic;
	signal   C440TRCBRANCHSTATUS_outdelay  :  std_logic_vector(0 to 2);
	signal   C440TRCCYCLE_outdelay  :  std_ulogic;
	signal   C440TRCEXECUTIONSTATUS_outdelay  :  std_logic_vector(0 to 4);
	signal   C440TRCTRACESTATUS_outdelay  :  std_logic_vector(0 to 6);
	signal   C440TRCTRIGGEREVENTOUT_outdelay  :  std_ulogic;
	signal   C440TRCTRIGGEREVENTTYPE_outdelay  :  std_logic_vector(0 to 13);
	signal   MIMCADDRESS_outdelay  :  std_logic_vector(0 to 35);
	signal   MIMCADDRESSVALID_outdelay  :  std_ulogic;
	signal   MIMCBANKCONFLICT_outdelay  :  std_ulogic;
	signal   MIMCBYTEENABLE_outdelay  :  std_logic_vector(0 to 15);
	signal   MIMCREADNOTWRITE_outdelay  :  std_ulogic;
	signal   MIMCROWCONFLICT_outdelay  :  std_ulogic;
	signal   MIMCWRITEDATA_outdelay  :  std_logic_vector(0 to 127);
	signal   MIMCWRITEDATAVALID_outdelay  :  std_ulogic;
	signal   PPCCPMINTERCONNECTBUSY_outdelay  :  std_ulogic;
	signal   PPCDSDCRACK_outdelay  :  std_ulogic;
	signal   PPCDSDCRTIMEOUTWAIT_outdelay  :  std_ulogic;
	signal   PPCDSDCRDBUSIN_outdelay  :  std_logic_vector(0 to 31);
	signal   PPCEICINTERCONNECTIRQ_outdelay  :  std_ulogic;

	signal   PLBPPCS0RNW_ipd  :  std_ulogic;
	signal   PLBPPCS1RNW_ipd  :  std_ulogic;
	signal   CPMDCRCLK_ipd  :  std_ulogic;
	signal   CPMDMA0LLCLK_ipd  :  std_ulogic;
	signal   CPMDMA1LLCLK_ipd  :  std_ulogic;
	signal   CPMDMA2LLCLK_ipd  :  std_ulogic;
	signal   CPMDMA3LLCLK_ipd  :  std_ulogic;
	signal   CPMINTERCONNECTCLKNTO1_ipd  :  std_ulogic;
	signal   CPMPPCMPLBCLK_ipd  :  std_ulogic;
	signal   CPMPPCS0PLBCLK_ipd  :  std_ulogic;
	signal   CPMPPCS1PLBCLK_ipd  :  std_ulogic;
	signal   DCRPPCDMACK_ipd  :  std_ulogic;
	signal   DCRPPCDMDBUSIN_ipd  :  std_logic_vector(0 to 31);
	signal   DCRPPCDMTIMEOUTWAIT_ipd  :  std_ulogic;
	signal   LLDMA0RSTENGINEREQ_ipd  :  std_ulogic;
	signal   LLDMA0RXD_ipd  :  std_logic_vector(0 to 31);
	signal   LLDMA0RXEOFN_ipd  :  std_ulogic;
	signal   LLDMA0RXEOPN_ipd  :  std_ulogic;
	signal   LLDMA0RXREM_ipd  :  std_logic_vector(0 to 3);
	signal   LLDMA0RXSOFN_ipd  :  std_ulogic;
	signal   LLDMA0RXSOPN_ipd  :  std_ulogic;
	signal   LLDMA0RXSRCRDYN_ipd  :  std_ulogic;
	signal   LLDMA0TXDSTRDYN_ipd  :  std_ulogic;
	signal   LLDMA1RSTENGINEREQ_ipd  :  std_ulogic;
	signal   LLDMA1RXD_ipd  :  std_logic_vector(0 to 31);
	signal   LLDMA1RXEOFN_ipd  :  std_ulogic;
	signal   LLDMA1RXEOPN_ipd  :  std_ulogic;
	signal   LLDMA1RXREM_ipd  :  std_logic_vector(0 to 3);
	signal   LLDMA1RXSOFN_ipd  :  std_ulogic;
	signal   LLDMA1RXSOPN_ipd  :  std_ulogic;
	signal   LLDMA1RXSRCRDYN_ipd  :  std_ulogic;
	signal   LLDMA1TXDSTRDYN_ipd  :  std_ulogic;
	signal   LLDMA2RSTENGINEREQ_ipd  :  std_ulogic;
	signal   LLDMA2RXD_ipd  :  std_logic_vector(0 to 31);
	signal   LLDMA2RXEOFN_ipd  :  std_ulogic;
	signal   LLDMA2RXEOPN_ipd  :  std_ulogic;
	signal   LLDMA2RXREM_ipd  :  std_logic_vector(0 to 3);
	signal   LLDMA2RXSOFN_ipd  :  std_ulogic;
	signal   LLDMA2RXSOPN_ipd  :  std_ulogic;
	signal   LLDMA2RXSRCRDYN_ipd  :  std_ulogic;
	signal   LLDMA2TXDSTRDYN_ipd  :  std_ulogic;
	signal   LLDMA3RSTENGINEREQ_ipd  :  std_ulogic;
	signal   LLDMA3RXD_ipd  :  std_logic_vector(0 to 31);
	signal   LLDMA3RXEOFN_ipd  :  std_ulogic;
	signal   LLDMA3RXEOPN_ipd  :  std_ulogic;
	signal   LLDMA3RXREM_ipd  :  std_logic_vector(0 to 3);
	signal   LLDMA3RXSOFN_ipd  :  std_ulogic;
	signal   LLDMA3RXSOPN_ipd  :  std_ulogic;
	signal   LLDMA3RXSRCRDYN_ipd  :  std_ulogic;
	signal   LLDMA3TXDSTRDYN_ipd  :  std_ulogic;
	signal   PLBPPCMADDRACK_ipd  :  std_ulogic;
	signal   PLBPPCMMBUSY_ipd  :  std_ulogic;
	signal   PLBPPCMMIRQ_ipd  :  std_ulogic;
	signal   PLBPPCMMRDERR_ipd  :  std_ulogic;
	signal   PLBPPCMMWRERR_ipd  :  std_ulogic;
	signal   PLBPPCMRDBTERM_ipd  :  std_ulogic;
	signal   PLBPPCMRDDACK_ipd  :  std_ulogic;
	signal   PLBPPCMRDDBUS_ipd  :  std_logic_vector(0 to 127);
	signal   PLBPPCMRDPENDPRI_ipd  :  std_logic_vector(0 to 1);
	signal   PLBPPCMRDPENDREQ_ipd  :  std_ulogic;
	signal   PLBPPCMRDWDADDR_ipd  :  std_logic_vector(0 to 3);
	signal   PLBPPCMREARBITRATE_ipd  :  std_ulogic;
	signal   PLBPPCMREQPRI_ipd  :  std_logic_vector(0 to 1);
	signal   PLBPPCMSSIZE_ipd  :  std_logic_vector(0 to 1);
	signal   PLBPPCMTIMEOUT_ipd  :  std_ulogic;
	signal   PLBPPCMWRBTERM_ipd  :  std_ulogic;
	signal   PLBPPCMWRDACK_ipd  :  std_ulogic;
	signal   PLBPPCMWRPENDPRI_ipd  :  std_logic_vector(0 to 1);
	signal   PLBPPCMWRPENDREQ_ipd  :  std_ulogic;
	signal   PLBPPCS0ABORT_ipd  :  std_ulogic;
	signal   PLBPPCS0ABUS_ipd  :  std_logic_vector(0 to 31);
	signal   PLBPPCS0BE_ipd  :  std_logic_vector(0 to 15);
	signal   PLBPPCS0BUSLOCK_ipd  :  std_ulogic;
	signal   PLBPPCS0LOCKERR_ipd  :  std_ulogic;
	signal   PLBPPCS0MASTERID_ipd  :  std_logic_vector(0 to 1);
	signal   PLBPPCS0MSIZE_ipd  :  std_logic_vector(0 to 1);
	signal   PLBPPCS0PAVALID_ipd  :  std_ulogic;
	signal   PLBPPCS0RDBURST_ipd  :  std_ulogic;
	signal   PLBPPCS0RDPENDPRI_ipd  :  std_logic_vector(0 to 1);
	signal   PLBPPCS0RDPENDREQ_ipd  :  std_ulogic;
	signal   PLBPPCS0RDPRIM_ipd  :  std_ulogic;
	signal   PLBPPCS0REQPRI_ipd  :  std_logic_vector(0 to 1);
	signal   PLBPPCS0SAVALID_ipd  :  std_ulogic;
	signal   PLBPPCS0SIZE_ipd  :  std_logic_vector(0 to 3);
	signal   PLBPPCS0TATTRIBUTE_ipd  :  std_logic_vector(0 to 15);
	signal   PLBPPCS0TYPE_ipd  :  std_logic_vector(0 to 2);
	signal   PLBPPCS0UABUS_ipd  :  std_logic_vector(28 to 31);
	signal   PLBPPCS0WRBURST_ipd  :  std_ulogic;
	signal   PLBPPCS0WRDBUS_ipd  :  std_logic_vector(0 to 127);
	signal   PLBPPCS0WRPENDPRI_ipd  :  std_logic_vector(0 to 1);
	signal   PLBPPCS0WRPENDREQ_ipd  :  std_ulogic;
	signal   PLBPPCS0WRPRIM_ipd  :  std_ulogic;
	signal   PLBPPCS1ABORT_ipd  :  std_ulogic;
	signal   PLBPPCS1ABUS_ipd  :  std_logic_vector(0 to 31);
	signal   PLBPPCS1BE_ipd  :  std_logic_vector(0 to 15);
	signal   PLBPPCS1BUSLOCK_ipd  :  std_ulogic;
	signal   PLBPPCS1LOCKERR_ipd  :  std_ulogic;
	signal   PLBPPCS1MASTERID_ipd  :  std_logic_vector(0 to 1);
	signal   PLBPPCS1MSIZE_ipd  :  std_logic_vector(0 to 1);
	signal   PLBPPCS1PAVALID_ipd  :  std_ulogic;
	signal   PLBPPCS1RDBURST_ipd  :  std_ulogic;
	signal   PLBPPCS1RDPENDPRI_ipd  :  std_logic_vector(0 to 1);
	signal   PLBPPCS1RDPENDREQ_ipd  :  std_ulogic;
	signal   PLBPPCS1RDPRIM_ipd  :  std_ulogic;
	signal   PLBPPCS1REQPRI_ipd  :  std_logic_vector(0 to 1);
	signal   PLBPPCS1SAVALID_ipd  :  std_ulogic;
	signal   PLBPPCS1SIZE_ipd  :  std_logic_vector(0 to 3);
	signal   PLBPPCS1TATTRIBUTE_ipd  :  std_logic_vector(0 to 15);
	signal   PLBPPCS1TYPE_ipd  :  std_logic_vector(0 to 2);
	signal   PLBPPCS1UABUS_ipd  :  std_logic_vector(28 to 31);
	signal   PLBPPCS1WRBURST_ipd  :  std_ulogic;
	signal   PLBPPCS1WRDBUS_ipd  :  std_logic_vector(0 to 127);
	signal   PLBPPCS1WRPENDPRI_ipd  :  std_logic_vector(0 to 1);
	signal   PLBPPCS1WRPENDREQ_ipd  :  std_ulogic;
	signal   PLBPPCS1WRPRIM_ipd  :  std_ulogic;
	signal   TIEDCRBASEADDR_ipd  :  std_logic_vector(0 to 1);
	signal   CPMC440CLK_ipd  :  std_ulogic;
	signal   CPMC440CLKEN_ipd  :  std_ulogic;
	signal   CPMC440CORECLOCKINACTIVE_ipd  :  std_ulogic;
	signal   CPMC440TIMERCLOCK_ipd  :  std_ulogic;
	signal   CPMFCMCLK_ipd  :  std_ulogic;
	signal   CPMINTERCONNECTCLK_ipd  :  std_ulogic;
	signal   CPMINTERCONNECTCLKEN_ipd  :  std_ulogic;
	signal   CPMMCCLK_ipd  :  std_ulogic;
	signal   DBGC440DEBUGHALT_ipd  :  std_ulogic;
	signal   DBGC440SYSTEMSTATUS_ipd  :  std_logic_vector(0 to 4);
	signal   DBGC440UNCONDDEBUGEVENT_ipd  :  std_ulogic;
	signal   DCRPPCDSABUS_ipd  :  std_logic_vector(0 to 9);
	signal   DCRPPCDSDBUSOUT_ipd  :  std_logic_vector(0 to 31);
	signal   DCRPPCDSREAD_ipd  :  std_ulogic;
	signal   DCRPPCDSWRITE_ipd  :  std_ulogic;
	signal   EICC440CRITIRQ_ipd  :  std_ulogic;
	signal   EICC440EXTIRQ_ipd  :  std_ulogic;
	signal   FCMAPUCONFIRMINSTR_ipd  :  std_ulogic;
	signal   FCMAPUCR_ipd  :  std_logic_vector(0 to 3);
	signal   FCMAPUDONE_ipd  :  std_ulogic;
	signal   FCMAPUEXCEPTION_ipd  :  std_ulogic;
	signal   FCMAPUFPSCRFEX_ipd  :  std_ulogic;
	signal   FCMAPURESULT_ipd  :  std_logic_vector(0 to 31);
	signal   FCMAPURESULTVALID_ipd  :  std_ulogic;
	signal   FCMAPUSLEEPNOTREADY_ipd  :  std_ulogic;
	signal   FCMAPUSTOREDATA_ipd  :  std_logic_vector(0 to 127);
	signal   JTGC440TCK_ipd  :  std_ulogic;
	signal   JTGC440TDI_ipd  :  std_ulogic;
	signal   JTGC440TMS_ipd  :  std_ulogic;
	signal   JTGC440TRSTNEG_ipd  :  std_ulogic;
	signal   MCMIADDRREADYTOACCEPT_ipd  :  std_ulogic;
	signal   MCMIREADDATA_ipd  :  std_logic_vector(0 to 127);
	signal   MCMIREADDATAERR_ipd  :  std_ulogic;
	signal   MCMIREADDATAVALID_ipd  :  std_ulogic;
	signal   RSTC440RESETCHIP_ipd  :  std_ulogic;
	signal   RSTC440RESETCORE_ipd  :  std_ulogic;
	signal   RSTC440RESETSYSTEM_ipd  :  std_ulogic;
	signal   TIEC440DCURDLDCACHEPLBPRIO_ipd  :  std_logic_vector(0 to 1);
	signal   TIEC440DCURDNONCACHEPLBPRIO_ipd  :  std_logic_vector(0 to 1);
	signal   TIEC440DCURDTOUCHPLBPRIO_ipd  :  std_logic_vector(0 to 1);
	signal   TIEC440DCURDURGENTPLBPRIO_ipd  :  std_logic_vector(0 to 1);
	signal   TIEC440DCUWRFLUSHPLBPRIO_ipd  :  std_logic_vector(0 to 1);
	signal   TIEC440DCUWRSTOREPLBPRIO_ipd  :  std_logic_vector(0 to 1);
	signal   TIEC440DCUWRURGENTPLBPRIO_ipd  :  std_logic_vector(0 to 1);
	signal   TIEC440ENDIANRESET_ipd  :  std_ulogic;
	signal   TIEC440ERPNRESET_ipd  :  std_logic_vector(0 to 3);
	signal   TIEC440ICURDFETCHPLBPRIO_ipd  :  std_logic_vector(0 to 1);
	signal   TIEC440ICURDSPECPLBPRIO_ipd  :  std_logic_vector(0 to 1);
	signal   TIEC440ICURDTOUCHPLBPRIO_ipd  :  std_logic_vector(0 to 1);
	signal   TIEC440PIR_ipd  :  std_logic_vector(28 to 31);
	signal   TIEC440PVR_ipd  :  std_logic_vector(28 to 31);
	signal   TIEC440USERRESET_ipd  :  std_logic_vector(0 to 3);
	signal   TRCC440TRACEDISABLE_ipd  :  std_ulogic;
	signal   TRCC440TRIGGEREVENTIN_ipd  :  std_ulogic;


	signal   PLBPPCS0RNW_indelay  :  std_ulogic;
	signal   PLBPPCS1RNW_indelay  :  std_ulogic;
	signal   CPMDCRCLK_indelay  :  std_ulogic;
	signal   CPMDMA0LLCLK_indelay  :  std_ulogic;
	signal   CPMDMA1LLCLK_indelay  :  std_ulogic;
	signal   CPMDMA2LLCLK_indelay  :  std_ulogic;
	signal   CPMDMA3LLCLK_indelay  :  std_ulogic;
	signal   CPMINTERCONNECTCLKNTO1_indelay  :  std_ulogic;
	signal   CPMPPCMPLBCLK_indelay  :  std_ulogic;
	signal   CPMPPCS0PLBCLK_indelay  :  std_ulogic;
	signal   CPMPPCS1PLBCLK_indelay  :  std_ulogic;
	signal   DCRPPCDMACK_indelay  :  std_ulogic;
	signal   DCRPPCDMDBUSIN_indelay  :  std_logic_vector(0 to 31);
	signal   DCRPPCDMTIMEOUTWAIT_indelay  :  std_ulogic;
	signal   LLDMA0RSTENGINEREQ_indelay  :  std_ulogic;
	signal   LLDMA0RXD_indelay  :  std_logic_vector(0 to 31);
	signal   LLDMA0RXEOFN_indelay  :  std_ulogic;
	signal   LLDMA0RXEOPN_indelay  :  std_ulogic;
	signal   LLDMA0RXREM_indelay  :  std_logic_vector(0 to 3);
	signal   LLDMA0RXSOFN_indelay  :  std_ulogic;
	signal   LLDMA0RXSOPN_indelay  :  std_ulogic;
	signal   LLDMA0RXSRCRDYN_indelay  :  std_ulogic;
	signal   LLDMA0TXDSTRDYN_indelay  :  std_ulogic;
	signal   LLDMA1RSTENGINEREQ_indelay  :  std_ulogic;
	signal   LLDMA1RXD_indelay  :  std_logic_vector(0 to 31);
	signal   LLDMA1RXEOFN_indelay  :  std_ulogic;
	signal   LLDMA1RXEOPN_indelay  :  std_ulogic;
	signal   LLDMA1RXREM_indelay  :  std_logic_vector(0 to 3);
	signal   LLDMA1RXSOFN_indelay  :  std_ulogic;
	signal   LLDMA1RXSOPN_indelay  :  std_ulogic;
	signal   LLDMA1RXSRCRDYN_indelay  :  std_ulogic;
	signal   LLDMA1TXDSTRDYN_indelay  :  std_ulogic;
	signal   LLDMA2RSTENGINEREQ_indelay  :  std_ulogic;
	signal   LLDMA2RXD_indelay  :  std_logic_vector(0 to 31);
	signal   LLDMA2RXEOFN_indelay  :  std_ulogic;
	signal   LLDMA2RXEOPN_indelay  :  std_ulogic;
	signal   LLDMA2RXREM_indelay  :  std_logic_vector(0 to 3);
	signal   LLDMA2RXSOFN_indelay  :  std_ulogic;
	signal   LLDMA2RXSOPN_indelay  :  std_ulogic;
	signal   LLDMA2RXSRCRDYN_indelay  :  std_ulogic;
	signal   LLDMA2TXDSTRDYN_indelay  :  std_ulogic;
	signal   LLDMA3RSTENGINEREQ_indelay  :  std_ulogic;
	signal   LLDMA3RXD_indelay  :  std_logic_vector(0 to 31);
	signal   LLDMA3RXEOFN_indelay  :  std_ulogic;
	signal   LLDMA3RXEOPN_indelay  :  std_ulogic;
	signal   LLDMA3RXREM_indelay  :  std_logic_vector(0 to 3);
	signal   LLDMA3RXSOFN_indelay  :  std_ulogic;
	signal   LLDMA3RXSOPN_indelay  :  std_ulogic;
	signal   LLDMA3RXSRCRDYN_indelay  :  std_ulogic;
	signal   LLDMA3TXDSTRDYN_indelay  :  std_ulogic;
	signal   PLBPPCMADDRACK_indelay  :  std_ulogic;
	signal   PLBPPCMMBUSY_indelay  :  std_ulogic;
	signal   PLBPPCMMIRQ_indelay  :  std_ulogic;
	signal   PLBPPCMMRDERR_indelay  :  std_ulogic;
	signal   PLBPPCMMWRERR_indelay  :  std_ulogic;
	signal   PLBPPCMRDBTERM_indelay  :  std_ulogic;
	signal   PLBPPCMRDDACK_indelay  :  std_ulogic;
	signal   PLBPPCMRDDBUS_indelay  :  std_logic_vector(0 to 127);
	signal   PLBPPCMRDPENDPRI_indelay  :  std_logic_vector(0 to 1);
	signal   PLBPPCMRDPENDREQ_indelay  :  std_ulogic;
	signal   PLBPPCMRDWDADDR_indelay  :  std_logic_vector(0 to 3);
	signal   PLBPPCMREARBITRATE_indelay  :  std_ulogic;
	signal   PLBPPCMREQPRI_indelay  :  std_logic_vector(0 to 1);
	signal   PLBPPCMSSIZE_indelay  :  std_logic_vector(0 to 1);
	signal   PLBPPCMTIMEOUT_indelay  :  std_ulogic;
	signal   PLBPPCMWRBTERM_indelay  :  std_ulogic;
	signal   PLBPPCMWRDACK_indelay  :  std_ulogic;
	signal   PLBPPCMWRPENDPRI_indelay  :  std_logic_vector(0 to 1);
	signal   PLBPPCMWRPENDREQ_indelay  :  std_ulogic;
	signal   PLBPPCS0ABORT_indelay  :  std_ulogic;
	signal   PLBPPCS0ABUS_indelay  :  std_logic_vector(0 to 31);
	signal   PLBPPCS0BE_indelay  :  std_logic_vector(0 to 15);
	signal   PLBPPCS0BUSLOCK_indelay  :  std_ulogic;
	signal   PLBPPCS0LOCKERR_indelay  :  std_ulogic;
	signal   PLBPPCS0MASTERID_indelay  :  std_logic_vector(0 to 1);
	signal   PLBPPCS0MSIZE_indelay  :  std_logic_vector(0 to 1);
	signal   PLBPPCS0PAVALID_indelay  :  std_ulogic;
	signal   PLBPPCS0RDBURST_indelay  :  std_ulogic;
	signal   PLBPPCS0RDPENDPRI_indelay  :  std_logic_vector(0 to 1);
	signal   PLBPPCS0RDPENDREQ_indelay  :  std_ulogic;
	signal   PLBPPCS0RDPRIM_indelay  :  std_ulogic;
	signal   PLBPPCS0REQPRI_indelay  :  std_logic_vector(0 to 1);
	signal   PLBPPCS0SAVALID_indelay  :  std_ulogic;
	signal   PLBPPCS0SIZE_indelay  :  std_logic_vector(0 to 3);
	signal   PLBPPCS0TATTRIBUTE_indelay  :  std_logic_vector(0 to 15);
	signal   PLBPPCS0TYPE_indelay  :  std_logic_vector(0 to 2);
	signal   PLBPPCS0UABUS_indelay  :  std_logic_vector(28 to 31);
	signal   PLBPPCS0WRBURST_indelay  :  std_ulogic;
	signal   PLBPPCS0WRDBUS_indelay  :  std_logic_vector(0 to 127);
	signal   PLBPPCS0WRPENDPRI_indelay  :  std_logic_vector(0 to 1);
	signal   PLBPPCS0WRPENDREQ_indelay  :  std_ulogic;
	signal   PLBPPCS0WRPRIM_indelay  :  std_ulogic;
	signal   PLBPPCS1ABORT_indelay  :  std_ulogic;
	signal   PLBPPCS1ABUS_indelay  :  std_logic_vector(0 to 31);
	signal   PLBPPCS1BE_indelay  :  std_logic_vector(0 to 15);
	signal   PLBPPCS1BUSLOCK_indelay  :  std_ulogic;
	signal   PLBPPCS1LOCKERR_indelay  :  std_ulogic;
	signal   PLBPPCS1MASTERID_indelay  :  std_logic_vector(0 to 1);
	signal   PLBPPCS1MSIZE_indelay  :  std_logic_vector(0 to 1);
	signal   PLBPPCS1PAVALID_indelay  :  std_ulogic;
	signal   PLBPPCS1RDBURST_indelay  :  std_ulogic;
	signal   PLBPPCS1RDPENDPRI_indelay  :  std_logic_vector(0 to 1);
	signal   PLBPPCS1RDPENDREQ_indelay  :  std_ulogic;
	signal   PLBPPCS1RDPRIM_indelay  :  std_ulogic;
	signal   PLBPPCS1REQPRI_indelay  :  std_logic_vector(0 to 1);
	signal   PLBPPCS1SAVALID_indelay  :  std_ulogic;
	signal   PLBPPCS1SIZE_indelay  :  std_logic_vector(0 to 3);
	signal   PLBPPCS1TATTRIBUTE_indelay  :  std_logic_vector(0 to 15);
	signal   PLBPPCS1TYPE_indelay  :  std_logic_vector(0 to 2);
	signal   PLBPPCS1UABUS_indelay  :  std_logic_vector(28 to 31);
	signal   PLBPPCS1WRBURST_indelay  :  std_ulogic;
	signal   PLBPPCS1WRDBUS_indelay  :  std_logic_vector(0 to 127);
	signal   PLBPPCS1WRPENDPRI_indelay  :  std_logic_vector(0 to 1);
	signal   PLBPPCS1WRPENDREQ_indelay  :  std_ulogic;
	signal   PLBPPCS1WRPRIM_indelay  :  std_ulogic;
	signal   TIEDCRBASEADDR_indelay  :  std_logic_vector(0 to 1);
	signal   CPMC440CLK_indelay  :  std_ulogic;
	signal   CPMC440CLKEN_indelay  :  std_ulogic;
	signal   CPMC440CORECLOCKINACTIVE_indelay  :  std_ulogic;
	signal   CPMC440TIMERCLOCK_indelay  :  std_ulogic;
	signal   CPMFCMCLK_indelay  :  std_ulogic;
	signal   CPMINTERCONNECTCLK_indelay  :  std_ulogic;
	signal   CPMINTERCONNECTCLKEN_indelay  :  std_ulogic;
	signal   CPMMCCLK_indelay  :  std_ulogic;
	signal   DBGC440DEBUGHALT_indelay  :  std_ulogic;
	signal   DBGC440SYSTEMSTATUS_indelay  :  std_logic_vector(0 to 4);
	signal   DBGC440UNCONDDEBUGEVENT_indelay  :  std_ulogic;
	signal   DCRPPCDSABUS_indelay  :  std_logic_vector(0 to 9);
	signal   DCRPPCDSDBUSOUT_indelay  :  std_logic_vector(0 to 31);
	signal   DCRPPCDSREAD_indelay  :  std_ulogic;
	signal   DCRPPCDSWRITE_indelay  :  std_ulogic;
	signal   EICC440CRITIRQ_indelay  :  std_ulogic;
	signal   EICC440EXTIRQ_indelay  :  std_ulogic;
	signal   FCMAPUCONFIRMINSTR_indelay  :  std_ulogic;
	signal   FCMAPUCR_indelay  :  std_logic_vector(0 to 3);
	signal   FCMAPUDONE_indelay  :  std_ulogic;
	signal   FCMAPUEXCEPTION_indelay  :  std_ulogic;
	signal   FCMAPUFPSCRFEX_indelay  :  std_ulogic;
	signal   FCMAPURESULT_indelay  :  std_logic_vector(0 to 31);
	signal   FCMAPURESULTVALID_indelay  :  std_ulogic;
	signal   FCMAPUSLEEPNOTREADY_indelay  :  std_ulogic;
	signal   FCMAPUSTOREDATA_indelay  :  std_logic_vector(0 to 127);
	signal   JTGC440TCK_indelay  :  std_ulogic;
	signal   JTGC440TDI_indelay  :  std_ulogic;
	signal   JTGC440TMS_indelay  :  std_ulogic;
	signal   JTGC440TRSTNEG_indelay  :  std_ulogic;
	signal   MCMIADDRREADYTOACCEPT_indelay  :  std_ulogic;
	signal   MCMIREADDATA_indelay  :  std_logic_vector(0 to 127);
	signal   MCMIREADDATAERR_indelay  :  std_ulogic;
	signal   MCMIREADDATAVALID_indelay  :  std_ulogic;
	signal   RSTC440RESETCHIP_indelay  :  std_ulogic;
	signal   RSTC440RESETCORE_indelay  :  std_ulogic;
	signal   RSTC440RESETSYSTEM_indelay  :  std_ulogic;
	signal   TIEC440DCURDLDCACHEPLBPRIO_indelay  :  std_logic_vector(0 to 1);
	signal   TIEC440DCURDNONCACHEPLBPRIO_indelay  :  std_logic_vector(0 to 1);
	signal   TIEC440DCURDTOUCHPLBPRIO_indelay  :  std_logic_vector(0 to 1);
	signal   TIEC440DCURDURGENTPLBPRIO_indelay  :  std_logic_vector(0 to 1);
	signal   TIEC440DCUWRFLUSHPLBPRIO_indelay  :  std_logic_vector(0 to 1);
	signal   TIEC440DCUWRSTOREPLBPRIO_indelay  :  std_logic_vector(0 to 1);
	signal   TIEC440DCUWRURGENTPLBPRIO_indelay  :  std_logic_vector(0 to 1);
	signal   TIEC440ENDIANRESET_indelay  :  std_ulogic;
	signal   TIEC440ERPNRESET_indelay  :  std_logic_vector(0 to 3);
	signal   TIEC440ICURDFETCHPLBPRIO_indelay  :  std_logic_vector(0 to 1);
	signal   TIEC440ICURDSPECPLBPRIO_indelay  :  std_logic_vector(0 to 1);
	signal   TIEC440ICURDTOUCHPLBPRIO_indelay  :  std_logic_vector(0 to 1);
	signal   TIEC440PIR_indelay  :  std_logic_vector(28 to 31);
	signal   TIEC440PVR_indelay  :  std_logic_vector(28 to 31);
	signal   TIEC440USERRESET_indelay  :  std_logic_vector(0 to 3);
	signal   TRCC440TRACEDISABLE_indelay  :  std_ulogic;
	signal   TRCC440TRIGGEREVENTIN_indelay  :  std_ulogic;

begin


	APUFCMDECFPUOP_out <= APUFCMDECFPUOP_outdelay after OUT_DELAY;
	APUFCMDECLDSTXFERSIZE_out <= APUFCMDECLDSTXFERSIZE_outdelay after OUT_DELAY;
	APUFCMDECLOAD_out <= APUFCMDECLOAD_outdelay after OUT_DELAY;
	APUFCMDECNONAUTON_out <= APUFCMDECNONAUTON_outdelay after OUT_DELAY;
	APUFCMDECSTORE_out <= APUFCMDECSTORE_outdelay after OUT_DELAY;
	APUFCMDECUDIVALID_out <= APUFCMDECUDIVALID_outdelay after OUT_DELAY;
	APUFCMDECUDI_out <= APUFCMDECUDI_outdelay after OUT_DELAY;
	APUFCMENDIAN_out <= APUFCMENDIAN_outdelay after OUT_DELAY;
	APUFCMFLUSH_out <= APUFCMFLUSH_outdelay after OUT_DELAY;
	APUFCMINSTRUCTION_out <= APUFCMINSTRUCTION_outdelay after OUT_DELAY;
	APUFCMINSTRVALID_out <= APUFCMINSTRVALID_outdelay after OUT_DELAY;
	APUFCMLOADBYTEADDR_out <= APUFCMLOADBYTEADDR_outdelay after OUT_DELAY;
	APUFCMLOADDATA_out <= APUFCMLOADDATA_outdelay after OUT_DELAY;
	APUFCMLOADDVALID_out <= APUFCMLOADDVALID_outdelay after OUT_DELAY;
	APUFCMMSRFE0_out <= APUFCMMSRFE0_outdelay after OUT_DELAY;
	APUFCMMSRFE1_out <= APUFCMMSRFE1_outdelay after OUT_DELAY;
	APUFCMNEXTINSTRREADY_out <= APUFCMNEXTINSTRREADY_outdelay after OUT_DELAY;
	APUFCMOPERANDVALID_out <= APUFCMOPERANDVALID_outdelay after OUT_DELAY;
	APUFCMRADATA_out <= APUFCMRADATA_outdelay after OUT_DELAY;
	APUFCMRBDATA_out <= APUFCMRBDATA_outdelay after OUT_DELAY;
	APUFCMWRITEBACKOK_out <= APUFCMWRITEBACKOK_outdelay after OUT_DELAY;
	C440CPMCORESLEEPREQ_out <= C440CPMCORESLEEPREQ_outdelay after OUT_DELAY;
	C440CPMDECIRPTREQ_out <= C440CPMDECIRPTREQ_outdelay after OUT_DELAY;
	C440CPMFITIRPTREQ_out <= C440CPMFITIRPTREQ_outdelay after OUT_DELAY;
	C440CPMMSRCE_out <= C440CPMMSRCE_outdelay after OUT_DELAY;
	C440CPMMSREE_out <= C440CPMMSREE_outdelay after OUT_DELAY;
	C440CPMTIMERRESETREQ_out <= C440CPMTIMERRESETREQ_outdelay after OUT_DELAY;
	C440CPMWDIRPTREQ_out <= C440CPMWDIRPTREQ_outdelay after OUT_DELAY;
	C440DBGSYSTEMCONTROL_out <= C440DBGSYSTEMCONTROL_outdelay after OUT_DELAY;
	C440JTGTDOEN_out <= C440JTGTDOEN_outdelay after OUT_DELAY;
	C440JTGTDO_out <= C440JTGTDO_outdelay after OUT_DELAY;
	C440MACHINECHECK_out <= C440MACHINECHECK_outdelay after OUT_DELAY;
	C440RSTCHIPRESETREQ_out <= C440RSTCHIPRESETREQ_outdelay after OUT_DELAY;
	C440RSTCORERESETREQ_out <= C440RSTCORERESETREQ_outdelay after OUT_DELAY;
	C440RSTSYSTEMRESETREQ_out <= C440RSTSYSTEMRESETREQ_outdelay after OUT_DELAY;
	C440TRCBRANCHSTATUS_out <= C440TRCBRANCHSTATUS_outdelay after OUT_DELAY;
	C440TRCCYCLE_out <= C440TRCCYCLE_outdelay after OUT_DELAY;
	C440TRCEXECUTIONSTATUS_out <= C440TRCEXECUTIONSTATUS_outdelay after OUT_DELAY;
	C440TRCTRACESTATUS_out <= C440TRCTRACESTATUS_outdelay after OUT_DELAY;
	C440TRCTRIGGEREVENTOUT_out <= C440TRCTRIGGEREVENTOUT_outdelay after OUT_DELAY;
	C440TRCTRIGGEREVENTTYPE_out <= C440TRCTRIGGEREVENTTYPE_outdelay after OUT_DELAY;
	DMA0LLRSTENGINEACK_out <= DMA0LLRSTENGINEACK_outdelay after OUT_DELAY;
	DMA0LLRXDSTRDYN_out <= DMA0LLRXDSTRDYN_outdelay after OUT_DELAY;
	DMA0LLTXD_out <= DMA0LLTXD_outdelay after OUT_DELAY;
	DMA0LLTXEOFN_out <= DMA0LLTXEOFN_outdelay after OUT_DELAY;
	DMA0LLTXEOPN_out <= DMA0LLTXEOPN_outdelay after OUT_DELAY;
	DMA0LLTXREM_out <= DMA0LLTXREM_outdelay after OUT_DELAY;
	DMA0LLTXSOFN_out <= DMA0LLTXSOFN_outdelay after OUT_DELAY;
	DMA0LLTXSOPN_out <= DMA0LLTXSOPN_outdelay after OUT_DELAY;
	DMA0LLTXSRCRDYN_out <= DMA0LLTXSRCRDYN_outdelay after OUT_DELAY;
	DMA0RXIRQ_out <= DMA0RXIRQ_outdelay after OUT_DELAY;
	DMA0TXIRQ_out <= DMA0TXIRQ_outdelay after OUT_DELAY;
	DMA1LLRSTENGINEACK_out <= DMA1LLRSTENGINEACK_outdelay after OUT_DELAY;
	DMA1LLRXDSTRDYN_out <= DMA1LLRXDSTRDYN_outdelay after OUT_DELAY;
	DMA1LLTXD_out <= DMA1LLTXD_outdelay after OUT_DELAY;
	DMA1LLTXEOFN_out <= DMA1LLTXEOFN_outdelay after OUT_DELAY;
	DMA1LLTXEOPN_out <= DMA1LLTXEOPN_outdelay after OUT_DELAY;
	DMA1LLTXREM_out <= DMA1LLTXREM_outdelay after OUT_DELAY;
	DMA1LLTXSOFN_out <= DMA1LLTXSOFN_outdelay after OUT_DELAY;
	DMA1LLTXSOPN_out <= DMA1LLTXSOPN_outdelay after OUT_DELAY;
	DMA1LLTXSRCRDYN_out <= DMA1LLTXSRCRDYN_outdelay after OUT_DELAY;
	DMA1RXIRQ_out <= DMA1RXIRQ_outdelay after OUT_DELAY;
	DMA1TXIRQ_out <= DMA1TXIRQ_outdelay after OUT_DELAY;
	DMA2LLRSTENGINEACK_out <= DMA2LLRSTENGINEACK_outdelay after OUT_DELAY;
	DMA2LLRXDSTRDYN_out <= DMA2LLRXDSTRDYN_outdelay after OUT_DELAY;
	DMA2LLTXD_out <= DMA2LLTXD_outdelay after OUT_DELAY;
	DMA2LLTXEOFN_out <= DMA2LLTXEOFN_outdelay after OUT_DELAY;
	DMA2LLTXEOPN_out <= DMA2LLTXEOPN_outdelay after OUT_DELAY;
	DMA2LLTXREM_out <= DMA2LLTXREM_outdelay after OUT_DELAY;
	DMA2LLTXSOFN_out <= DMA2LLTXSOFN_outdelay after OUT_DELAY;
	DMA2LLTXSOPN_out <= DMA2LLTXSOPN_outdelay after OUT_DELAY;
	DMA2LLTXSRCRDYN_out <= DMA2LLTXSRCRDYN_outdelay after OUT_DELAY;
	DMA2RXIRQ_out <= DMA2RXIRQ_outdelay after OUT_DELAY;
	DMA2TXIRQ_out <= DMA2TXIRQ_outdelay after OUT_DELAY;
	DMA3LLRSTENGINEACK_out <= DMA3LLRSTENGINEACK_outdelay after OUT_DELAY;
	DMA3LLRXDSTRDYN_out <= DMA3LLRXDSTRDYN_outdelay after OUT_DELAY;
	DMA3LLTXD_out <= DMA3LLTXD_outdelay after OUT_DELAY;
	DMA3LLTXEOFN_out <= DMA3LLTXEOFN_outdelay after OUT_DELAY;
	DMA3LLTXEOPN_out <= DMA3LLTXEOPN_outdelay after OUT_DELAY;
	DMA3LLTXREM_out <= DMA3LLTXREM_outdelay after OUT_DELAY;
	DMA3LLTXSOFN_out <= DMA3LLTXSOFN_outdelay after OUT_DELAY;
	DMA3LLTXSOPN_out <= DMA3LLTXSOPN_outdelay after OUT_DELAY;
	DMA3LLTXSRCRDYN_out <= DMA3LLTXSRCRDYN_outdelay after OUT_DELAY;
	DMA3RXIRQ_out <= DMA3RXIRQ_outdelay after OUT_DELAY;
	DMA3TXIRQ_out <= DMA3TXIRQ_outdelay after OUT_DELAY;
	MIMCADDRESSVALID_out <= MIMCADDRESSVALID_outdelay after OUT_DELAY;
	MIMCADDRESS_out <= MIMCADDRESS_outdelay after OUT_DELAY;
	MIMCBANKCONFLICT_out <= MIMCBANKCONFLICT_outdelay after OUT_DELAY;
	MIMCBYTEENABLE_out <= MIMCBYTEENABLE_outdelay after OUT_DELAY;
	MIMCREADNOTWRITE_out <= MIMCREADNOTWRITE_outdelay after OUT_DELAY;
	MIMCROWCONFLICT_out <= MIMCROWCONFLICT_outdelay after OUT_DELAY;
	MIMCWRITEDATAVALID_out <= MIMCWRITEDATAVALID_outdelay after OUT_DELAY;
	MIMCWRITEDATA_out <= MIMCWRITEDATA_outdelay after OUT_DELAY;
	PPCCPMINTERCONNECTBUSY_out <= PPCCPMINTERCONNECTBUSY_outdelay after OUT_DELAY;
	PPCDMDCRABUS_out <= PPCDMDCRABUS_outdelay after OUT_DELAY;
	PPCDMDCRDBUSOUT_out <= PPCDMDCRDBUSOUT_outdelay after OUT_DELAY;
	PPCDMDCRREAD_out <= PPCDMDCRREAD_outdelay after OUT_DELAY;
	PPCDMDCRUABUS_out <= PPCDMDCRUABUS_outdelay after OUT_DELAY;
	PPCDMDCRWRITE_out <= PPCDMDCRWRITE_outdelay after OUT_DELAY;
	PPCDSDCRACK_out <= PPCDSDCRACK_outdelay after OUT_DELAY;
	PPCDSDCRDBUSIN_out <= PPCDSDCRDBUSIN_outdelay after OUT_DELAY;
	PPCDSDCRTIMEOUTWAIT_out <= PPCDSDCRTIMEOUTWAIT_outdelay after OUT_DELAY;
	PPCEICINTERCONNECTIRQ_out <= PPCEICINTERCONNECTIRQ_outdelay after OUT_DELAY;
	PPCMPLBABORT_out <= PPCMPLBABORT_outdelay after OUT_DELAY;
	PPCMPLBABUS_out <= PPCMPLBABUS_outdelay after OUT_DELAY;
	PPCMPLBBE_out <= PPCMPLBBE_outdelay after OUT_DELAY;
	PPCMPLBBUSLOCK_out <= PPCMPLBBUSLOCK_outdelay after OUT_DELAY;
	PPCMPLBLOCKERR_out <= PPCMPLBLOCKERR_outdelay after OUT_DELAY;
	PPCMPLBPRIORITY_out <= PPCMPLBPRIORITY_outdelay after OUT_DELAY;
	PPCMPLBRDBURST_out <= PPCMPLBRDBURST_outdelay after OUT_DELAY;
	PPCMPLBREQUEST_out <= PPCMPLBREQUEST_outdelay after OUT_DELAY;
	PPCMPLBRNW_out <= PPCMPLBRNW_outdelay after OUT_DELAY;
	PPCMPLBSIZE_out <= PPCMPLBSIZE_outdelay after OUT_DELAY;
	PPCMPLBTATTRIBUTE_out <= PPCMPLBTATTRIBUTE_outdelay after OUT_DELAY;
	PPCMPLBTYPE_out <= PPCMPLBTYPE_outdelay after OUT_DELAY;
	PPCMPLBUABUS_out <= PPCMPLBUABUS_outdelay after OUT_DELAY;
	PPCMPLBWRBURST_out <= PPCMPLBWRBURST_outdelay after OUT_DELAY;
	PPCMPLBWRDBUS_out <= PPCMPLBWRDBUS_outdelay after OUT_DELAY;
	PPCS0PLBADDRACK_out <= PPCS0PLBADDRACK_outdelay after OUT_DELAY;
	PPCS0PLBMBUSY_out <= PPCS0PLBMBUSY_outdelay after OUT_DELAY;
	PPCS0PLBMIRQ_out <= PPCS0PLBMIRQ_outdelay after OUT_DELAY;
	PPCS0PLBMRDERR_out <= PPCS0PLBMRDERR_outdelay after OUT_DELAY;
	PPCS0PLBMWRERR_out <= PPCS0PLBMWRERR_outdelay after OUT_DELAY;
	PPCS0PLBRDBTERM_out <= PPCS0PLBRDBTERM_outdelay after OUT_DELAY;
	PPCS0PLBRDCOMP_out <= PPCS0PLBRDCOMP_outdelay after OUT_DELAY;
	PPCS0PLBRDDACK_out <= PPCS0PLBRDDACK_outdelay after OUT_DELAY;
	PPCS0PLBRDDBUS_out <= PPCS0PLBRDDBUS_outdelay after OUT_DELAY;
	PPCS0PLBRDWDADDR_out <= PPCS0PLBRDWDADDR_outdelay after OUT_DELAY;
	PPCS0PLBREARBITRATE_out <= PPCS0PLBREARBITRATE_outdelay after OUT_DELAY;
	PPCS0PLBSSIZE_out <= PPCS0PLBSSIZE_outdelay after OUT_DELAY;
	PPCS0PLBWAIT_out <= PPCS0PLBWAIT_outdelay after OUT_DELAY;
	PPCS0PLBWRBTERM_out <= PPCS0PLBWRBTERM_outdelay after OUT_DELAY;
	PPCS0PLBWRCOMP_out <= PPCS0PLBWRCOMP_outdelay after OUT_DELAY;
	PPCS0PLBWRDACK_out <= PPCS0PLBWRDACK_outdelay after OUT_DELAY;
	PPCS1PLBADDRACK_out <= PPCS1PLBADDRACK_outdelay after OUT_DELAY;
	PPCS1PLBMBUSY_out <= PPCS1PLBMBUSY_outdelay after OUT_DELAY;
	PPCS1PLBMIRQ_out <= PPCS1PLBMIRQ_outdelay after OUT_DELAY;
	PPCS1PLBMRDERR_out <= PPCS1PLBMRDERR_outdelay after OUT_DELAY;
	PPCS1PLBMWRERR_out <= PPCS1PLBMWRERR_outdelay after OUT_DELAY;
	PPCS1PLBRDBTERM_out <= PPCS1PLBRDBTERM_outdelay after OUT_DELAY;
	PPCS1PLBRDCOMP_out <= PPCS1PLBRDCOMP_outdelay after OUT_DELAY;
	PPCS1PLBRDDACK_out <= PPCS1PLBRDDACK_outdelay after OUT_DELAY;
	PPCS1PLBRDDBUS_out <= PPCS1PLBRDDBUS_outdelay after OUT_DELAY;
	PPCS1PLBRDWDADDR_out <= PPCS1PLBRDWDADDR_outdelay after OUT_DELAY;
	PPCS1PLBREARBITRATE_out <= PPCS1PLBREARBITRATE_outdelay after OUT_DELAY;
	PPCS1PLBSSIZE_out <= PPCS1PLBSSIZE_outdelay after OUT_DELAY;
	PPCS1PLBWAIT_out <= PPCS1PLBWAIT_outdelay after OUT_DELAY;
	PPCS1PLBWRBTERM_out <= PPCS1PLBWRBTERM_outdelay after OUT_DELAY;
	PPCS1PLBWRCOMP_out <= PPCS1PLBWRCOMP_outdelay after OUT_DELAY;
	PPCS1PLBWRDACK_out <= PPCS1PLBWRDACK_outdelay after OUT_DELAY;

	CPMC440CLK_ipd <= CPMC440CLK after ZERO_DELAY;
	CPMC440TIMERCLOCK_ipd <= CPMC440TIMERCLOCK after ZERO_DELAY;
	CPMDCRCLK_ipd <= CPMDCRCLK after ZERO_DELAY;
	CPMDMA0LLCLK_ipd <= CPMDMA0LLCLK after ZERO_DELAY;
	CPMDMA1LLCLK_ipd <= CPMDMA1LLCLK after ZERO_DELAY;
	CPMDMA2LLCLK_ipd <= CPMDMA2LLCLK after ZERO_DELAY;
	CPMDMA3LLCLK_ipd <= CPMDMA3LLCLK after ZERO_DELAY;
	CPMFCMCLK_ipd <= CPMFCMCLK after ZERO_DELAY;
	CPMINTERCONNECTCLK_ipd <= CPMINTERCONNECTCLK after ZERO_DELAY;
	CPMMCCLK_ipd <= CPMMCCLK after ZERO_DELAY;
	CPMPPCMPLBCLK_ipd <= CPMPPCMPLBCLK after ZERO_DELAY;
	CPMPPCS0PLBCLK_ipd <= CPMPPCS0PLBCLK after ZERO_DELAY;
	CPMPPCS1PLBCLK_ipd <= CPMPPCS1PLBCLK after ZERO_DELAY;
	JTGC440TCK_ipd <= JTGC440TCK after ZERO_DELAY;

	CPMC440CLKEN_ipd <= CPMC440CLKEN after ZERO_DELAY;
	CPMC440CORECLOCKINACTIVE_ipd <= CPMC440CORECLOCKINACTIVE after ZERO_DELAY;
	CPMINTERCONNECTCLKEN_ipd <= CPMINTERCONNECTCLKEN after ZERO_DELAY;
	CPMINTERCONNECTCLKNTO1_ipd <= CPMINTERCONNECTCLKNTO1 after ZERO_DELAY;
	DBGC440DEBUGHALT_ipd <= DBGC440DEBUGHALT after ZERO_DELAY;
	DBGC440SYSTEMSTATUS_ipd <= DBGC440SYSTEMSTATUS after ZERO_DELAY;
	DBGC440UNCONDDEBUGEVENT_ipd <= DBGC440UNCONDDEBUGEVENT after ZERO_DELAY;
	DCRPPCDMACK_ipd <= DCRPPCDMACK after ZERO_DELAY;
	DCRPPCDMDBUSIN_ipd <= DCRPPCDMDBUSIN after ZERO_DELAY;
	DCRPPCDMTIMEOUTWAIT_ipd <= DCRPPCDMTIMEOUTWAIT after ZERO_DELAY;
	DCRPPCDSABUS_ipd <= DCRPPCDSABUS after ZERO_DELAY;
	DCRPPCDSDBUSOUT_ipd <= DCRPPCDSDBUSOUT after ZERO_DELAY;
	DCRPPCDSREAD_ipd <= DCRPPCDSREAD after ZERO_DELAY;
	DCRPPCDSWRITE_ipd <= DCRPPCDSWRITE after ZERO_DELAY;
	EICC440CRITIRQ_ipd <= EICC440CRITIRQ after ZERO_DELAY;
	EICC440EXTIRQ_ipd <= EICC440EXTIRQ after ZERO_DELAY;
	FCMAPUCONFIRMINSTR_ipd <= FCMAPUCONFIRMINSTR after ZERO_DELAY;
	FCMAPUCR_ipd <= FCMAPUCR after ZERO_DELAY;
	FCMAPUDONE_ipd <= FCMAPUDONE after ZERO_DELAY;
	FCMAPUEXCEPTION_ipd <= FCMAPUEXCEPTION after ZERO_DELAY;
	FCMAPUFPSCRFEX_ipd <= FCMAPUFPSCRFEX after ZERO_DELAY;
	FCMAPURESULTVALID_ipd <= FCMAPURESULTVALID after ZERO_DELAY;
	FCMAPURESULT_ipd <= FCMAPURESULT after ZERO_DELAY;
	FCMAPUSLEEPNOTREADY_ipd <= FCMAPUSLEEPNOTREADY after ZERO_DELAY;
	FCMAPUSTOREDATA_ipd <= FCMAPUSTOREDATA after ZERO_DELAY;
	JTGC440TDI_ipd <= JTGC440TDI after ZERO_DELAY;
	JTGC440TMS_ipd <= JTGC440TMS after ZERO_DELAY;
	JTGC440TRSTNEG_ipd <= JTGC440TRSTNEG after ZERO_DELAY;
	LLDMA0RSTENGINEREQ_ipd <= LLDMA0RSTENGINEREQ after ZERO_DELAY;
	LLDMA0RXD_ipd <= LLDMA0RXD after ZERO_DELAY;
	LLDMA0RXEOFN_ipd <= LLDMA0RXEOFN after ZERO_DELAY;
	LLDMA0RXEOPN_ipd <= LLDMA0RXEOPN after ZERO_DELAY;
	LLDMA0RXREM_ipd <= LLDMA0RXREM after ZERO_DELAY;
	LLDMA0RXSOFN_ipd <= LLDMA0RXSOFN after ZERO_DELAY;
	LLDMA0RXSOPN_ipd <= LLDMA0RXSOPN after ZERO_DELAY;
	LLDMA0RXSRCRDYN_ipd <= LLDMA0RXSRCRDYN after ZERO_DELAY;
	LLDMA0TXDSTRDYN_ipd <= LLDMA0TXDSTRDYN after ZERO_DELAY;
	LLDMA1RSTENGINEREQ_ipd <= LLDMA1RSTENGINEREQ after ZERO_DELAY;
	LLDMA1RXD_ipd <= LLDMA1RXD after ZERO_DELAY;
	LLDMA1RXEOFN_ipd <= LLDMA1RXEOFN after ZERO_DELAY;
	LLDMA1RXEOPN_ipd <= LLDMA1RXEOPN after ZERO_DELAY;
	LLDMA1RXREM_ipd <= LLDMA1RXREM after ZERO_DELAY;
	LLDMA1RXSOFN_ipd <= LLDMA1RXSOFN after ZERO_DELAY;
	LLDMA1RXSOPN_ipd <= LLDMA1RXSOPN after ZERO_DELAY;
	LLDMA1RXSRCRDYN_ipd <= LLDMA1RXSRCRDYN after ZERO_DELAY;
	LLDMA1TXDSTRDYN_ipd <= LLDMA1TXDSTRDYN after ZERO_DELAY;
	LLDMA2RSTENGINEREQ_ipd <= LLDMA2RSTENGINEREQ after ZERO_DELAY;
	LLDMA2RXD_ipd <= LLDMA2RXD after ZERO_DELAY;
	LLDMA2RXEOFN_ipd <= LLDMA2RXEOFN after ZERO_DELAY;
	LLDMA2RXEOPN_ipd <= LLDMA2RXEOPN after ZERO_DELAY;
	LLDMA2RXREM_ipd <= LLDMA2RXREM after ZERO_DELAY;
	LLDMA2RXSOFN_ipd <= LLDMA2RXSOFN after ZERO_DELAY;
	LLDMA2RXSOPN_ipd <= LLDMA2RXSOPN after ZERO_DELAY;
	LLDMA2RXSRCRDYN_ipd <= LLDMA2RXSRCRDYN after ZERO_DELAY;
	LLDMA2TXDSTRDYN_ipd <= LLDMA2TXDSTRDYN after ZERO_DELAY;
	LLDMA3RSTENGINEREQ_ipd <= LLDMA3RSTENGINEREQ after ZERO_DELAY;
	LLDMA3RXD_ipd <= LLDMA3RXD after ZERO_DELAY;
	LLDMA3RXEOFN_ipd <= LLDMA3RXEOFN after ZERO_DELAY;
	LLDMA3RXEOPN_ipd <= LLDMA3RXEOPN after ZERO_DELAY;
	LLDMA3RXREM_ipd <= LLDMA3RXREM after ZERO_DELAY;
	LLDMA3RXSOFN_ipd <= LLDMA3RXSOFN after ZERO_DELAY;
	LLDMA3RXSOPN_ipd <= LLDMA3RXSOPN after ZERO_DELAY;
	LLDMA3RXSRCRDYN_ipd <= LLDMA3RXSRCRDYN after ZERO_DELAY;
	LLDMA3TXDSTRDYN_ipd <= LLDMA3TXDSTRDYN after ZERO_DELAY;
	MCMIADDRREADYTOACCEPT_ipd <= MCMIADDRREADYTOACCEPT after ZERO_DELAY;
	MCMIREADDATAERR_ipd <= MCMIREADDATAERR after ZERO_DELAY;
	MCMIREADDATAVALID_ipd <= MCMIREADDATAVALID after ZERO_DELAY;
	MCMIREADDATA_ipd <= MCMIREADDATA after ZERO_DELAY;
	PLBPPCMADDRACK_ipd <= PLBPPCMADDRACK after ZERO_DELAY;
	PLBPPCMMBUSY_ipd <= PLBPPCMMBUSY after ZERO_DELAY;
	PLBPPCMMIRQ_ipd <= PLBPPCMMIRQ after ZERO_DELAY;
	PLBPPCMMRDERR_ipd <= PLBPPCMMRDERR after ZERO_DELAY;
	PLBPPCMMWRERR_ipd <= PLBPPCMMWRERR after ZERO_DELAY;
	PLBPPCMRDBTERM_ipd <= PLBPPCMRDBTERM after ZERO_DELAY;
	PLBPPCMRDDACK_ipd <= PLBPPCMRDDACK after ZERO_DELAY;
	PLBPPCMRDDBUS_ipd <= PLBPPCMRDDBUS after ZERO_DELAY;
	PLBPPCMRDPENDPRI_ipd <= PLBPPCMRDPENDPRI after ZERO_DELAY;
	PLBPPCMRDPENDREQ_ipd <= PLBPPCMRDPENDREQ after ZERO_DELAY;
	PLBPPCMRDWDADDR_ipd <= PLBPPCMRDWDADDR after ZERO_DELAY;
	PLBPPCMREARBITRATE_ipd <= PLBPPCMREARBITRATE after ZERO_DELAY;
	PLBPPCMREQPRI_ipd <= PLBPPCMREQPRI after ZERO_DELAY;
	PLBPPCMSSIZE_ipd <= PLBPPCMSSIZE after ZERO_DELAY;
	PLBPPCMTIMEOUT_ipd <= PLBPPCMTIMEOUT after ZERO_DELAY;
	PLBPPCMWRBTERM_ipd <= PLBPPCMWRBTERM after ZERO_DELAY;
	PLBPPCMWRDACK_ipd <= PLBPPCMWRDACK after ZERO_DELAY;
	PLBPPCMWRPENDPRI_ipd <= PLBPPCMWRPENDPRI after ZERO_DELAY;
	PLBPPCMWRPENDREQ_ipd <= PLBPPCMWRPENDREQ after ZERO_DELAY;
	PLBPPCS0ABORT_ipd <= PLBPPCS0ABORT after ZERO_DELAY;
	PLBPPCS0ABUS_ipd <= PLBPPCS0ABUS after ZERO_DELAY;
	PLBPPCS0BE_ipd <= PLBPPCS0BE after ZERO_DELAY;
	PLBPPCS0BUSLOCK_ipd <= PLBPPCS0BUSLOCK after ZERO_DELAY;
	PLBPPCS0LOCKERR_ipd <= PLBPPCS0LOCKERR after ZERO_DELAY;
	PLBPPCS0MASTERID_ipd <= PLBPPCS0MASTERID after ZERO_DELAY;
	PLBPPCS0MSIZE_ipd <= PLBPPCS0MSIZE after ZERO_DELAY;
	PLBPPCS0PAVALID_ipd <= PLBPPCS0PAVALID after ZERO_DELAY;
	PLBPPCS0RDBURST_ipd <= PLBPPCS0RDBURST after ZERO_DELAY;
	PLBPPCS0RDPENDPRI_ipd <= PLBPPCS0RDPENDPRI after ZERO_DELAY;
	PLBPPCS0RDPENDREQ_ipd <= PLBPPCS0RDPENDREQ after ZERO_DELAY;
	PLBPPCS0RDPRIM_ipd <= PLBPPCS0RDPRIM after ZERO_DELAY;
	PLBPPCS0REQPRI_ipd <= PLBPPCS0REQPRI after ZERO_DELAY;
	PLBPPCS0RNW_ipd <= PLBPPCS0RNW after ZERO_DELAY;
	PLBPPCS0SAVALID_ipd <= PLBPPCS0SAVALID after ZERO_DELAY;
	PLBPPCS0SIZE_ipd <= PLBPPCS0SIZE after ZERO_DELAY;
	PLBPPCS0TATTRIBUTE_ipd <= PLBPPCS0TATTRIBUTE after ZERO_DELAY;
	PLBPPCS0TYPE_ipd <= PLBPPCS0TYPE after ZERO_DELAY;
	PLBPPCS0UABUS_ipd <= PLBPPCS0UABUS after ZERO_DELAY;
	PLBPPCS0WRBURST_ipd <= PLBPPCS0WRBURST after ZERO_DELAY;
	PLBPPCS0WRDBUS_ipd <= PLBPPCS0WRDBUS after ZERO_DELAY;
	PLBPPCS0WRPENDPRI_ipd <= PLBPPCS0WRPENDPRI after ZERO_DELAY;
	PLBPPCS0WRPENDREQ_ipd <= PLBPPCS0WRPENDREQ after ZERO_DELAY;
	PLBPPCS0WRPRIM_ipd <= PLBPPCS0WRPRIM after ZERO_DELAY;
	PLBPPCS1ABORT_ipd <= PLBPPCS1ABORT after ZERO_DELAY;
	PLBPPCS1ABUS_ipd <= PLBPPCS1ABUS after ZERO_DELAY;
	PLBPPCS1BE_ipd <= PLBPPCS1BE after ZERO_DELAY;
	PLBPPCS1BUSLOCK_ipd <= PLBPPCS1BUSLOCK after ZERO_DELAY;
	PLBPPCS1LOCKERR_ipd <= PLBPPCS1LOCKERR after ZERO_DELAY;
	PLBPPCS1MASTERID_ipd <= PLBPPCS1MASTERID after ZERO_DELAY;
	PLBPPCS1MSIZE_ipd <= PLBPPCS1MSIZE after ZERO_DELAY;
	PLBPPCS1PAVALID_ipd <= PLBPPCS1PAVALID after ZERO_DELAY;
	PLBPPCS1RDBURST_ipd <= PLBPPCS1RDBURST after ZERO_DELAY;
	PLBPPCS1RDPENDPRI_ipd <= PLBPPCS1RDPENDPRI after ZERO_DELAY;
	PLBPPCS1RDPENDREQ_ipd <= PLBPPCS1RDPENDREQ after ZERO_DELAY;
	PLBPPCS1RDPRIM_ipd <= PLBPPCS1RDPRIM after ZERO_DELAY;
	PLBPPCS1REQPRI_ipd <= PLBPPCS1REQPRI after ZERO_DELAY;
	PLBPPCS1RNW_ipd <= PLBPPCS1RNW after ZERO_DELAY;
	PLBPPCS1SAVALID_ipd <= PLBPPCS1SAVALID after ZERO_DELAY;
	PLBPPCS1SIZE_ipd <= PLBPPCS1SIZE after ZERO_DELAY;
	PLBPPCS1TATTRIBUTE_ipd <= PLBPPCS1TATTRIBUTE after ZERO_DELAY;
	PLBPPCS1TYPE_ipd <= PLBPPCS1TYPE after ZERO_DELAY;
	PLBPPCS1UABUS_ipd <= PLBPPCS1UABUS after ZERO_DELAY;
	PLBPPCS1WRBURST_ipd <= PLBPPCS1WRBURST after ZERO_DELAY;
	PLBPPCS1WRDBUS_ipd <= PLBPPCS1WRDBUS after ZERO_DELAY;
	PLBPPCS1WRPENDPRI_ipd <= PLBPPCS1WRPENDPRI after ZERO_DELAY;
	PLBPPCS1WRPENDREQ_ipd <= PLBPPCS1WRPENDREQ after ZERO_DELAY;
	PLBPPCS1WRPRIM_ipd <= PLBPPCS1WRPRIM after ZERO_DELAY;
	RSTC440RESETCHIP_ipd <= RSTC440RESETCHIP after ZERO_DELAY;
	RSTC440RESETCORE_ipd <= RSTC440RESETCORE after ZERO_DELAY;
	RSTC440RESETSYSTEM_ipd <= RSTC440RESETSYSTEM after ZERO_DELAY;
	TIEC440DCURDLDCACHEPLBPRIO_ipd <= TIEC440DCURDLDCACHEPLBPRIO after ZERO_DELAY;
	TIEC440DCURDNONCACHEPLBPRIO_ipd <= TIEC440DCURDNONCACHEPLBPRIO after ZERO_DELAY;
	TIEC440DCURDTOUCHPLBPRIO_ipd <= TIEC440DCURDTOUCHPLBPRIO after ZERO_DELAY;
	TIEC440DCURDURGENTPLBPRIO_ipd <= TIEC440DCURDURGENTPLBPRIO after ZERO_DELAY;
	TIEC440DCUWRFLUSHPLBPRIO_ipd <= TIEC440DCUWRFLUSHPLBPRIO after ZERO_DELAY;
	TIEC440DCUWRSTOREPLBPRIO_ipd <= TIEC440DCUWRSTOREPLBPRIO after ZERO_DELAY;
	TIEC440DCUWRURGENTPLBPRIO_ipd <= TIEC440DCUWRURGENTPLBPRIO after ZERO_DELAY;
	TIEC440ENDIANRESET_ipd <= TIEC440ENDIANRESET after ZERO_DELAY;
	TIEC440ERPNRESET_ipd <= TIEC440ERPNRESET after ZERO_DELAY;
	TIEC440ICURDFETCHPLBPRIO_ipd <= TIEC440ICURDFETCHPLBPRIO after ZERO_DELAY;
	TIEC440ICURDSPECPLBPRIO_ipd <= TIEC440ICURDSPECPLBPRIO after ZERO_DELAY;
	TIEC440ICURDTOUCHPLBPRIO_ipd <= TIEC440ICURDTOUCHPLBPRIO after ZERO_DELAY;
	TIEC440PIR_ipd <= TIEC440PIR after ZERO_DELAY;
	TIEC440PVR_ipd <= TIEC440PVR after ZERO_DELAY;
	TIEC440USERRESET_ipd <= TIEC440USERRESET after ZERO_DELAY;
	TIEDCRBASEADDR_ipd <= TIEDCRBASEADDR after ZERO_DELAY;
	TRCC440TRACEDISABLE_ipd <= TRCC440TRACEDISABLE after ZERO_DELAY;
	TRCC440TRIGGEREVENTIN_ipd <= TRCC440TRIGGEREVENTIN after ZERO_DELAY;


	CPMC440CLK_indelay <= CPMC440CLK_ipd after CLK_DELAY;
	CPMC440TIMERCLOCK_indelay <= CPMC440TIMERCLOCK_ipd after CLK_DELAY;
	CPMDCRCLK_indelay <= CPMDCRCLK_ipd after CLK_DELAY;
	CPMDMA0LLCLK_indelay <= CPMDMA0LLCLK_ipd after CLK_DELAY;
	CPMDMA1LLCLK_indelay <= CPMDMA1LLCLK_ipd after CLK_DELAY;
	CPMDMA2LLCLK_indelay <= CPMDMA2LLCLK_ipd after CLK_DELAY;
	CPMDMA3LLCLK_indelay <= CPMDMA3LLCLK_ipd after CLK_DELAY;
	CPMFCMCLK_indelay <= CPMFCMCLK_ipd after CLK_DELAY;
	CPMINTERCONNECTCLK_indelay <= CPMINTERCONNECTCLK_ipd after CLK_DELAY;
	CPMMCCLK_indelay <= CPMMCCLK_ipd after CLK_DELAY;
	CPMPPCMPLBCLK_indelay <= CPMPPCMPLBCLK_ipd after CLK_DELAY;
	CPMPPCS0PLBCLK_indelay <= CPMPPCS0PLBCLK_ipd after CLK_DELAY;
	CPMPPCS1PLBCLK_indelay <= CPMPPCS1PLBCLK_ipd after CLK_DELAY;
	JTGC440TCK_indelay <= JTGC440TCK_ipd after CLK_DELAY;

	CPMC440CLKEN_indelay <= CPMC440CLKEN_ipd after IN_DELAY;
	CPMC440CORECLOCKINACTIVE_indelay <= CPMC440CORECLOCKINACTIVE_ipd after IN_DELAY;
	CPMINTERCONNECTCLKEN_indelay <= CPMINTERCONNECTCLKEN_ipd after IN_DELAY;
	CPMINTERCONNECTCLKNTO1_indelay <= CPMINTERCONNECTCLKNTO1_ipd after IN_DELAY;
	DBGC440DEBUGHALT_indelay <= DBGC440DEBUGHALT_ipd after IN_DELAY;
	DBGC440SYSTEMSTATUS_indelay <= DBGC440SYSTEMSTATUS_ipd after IN_DELAY;
	DBGC440UNCONDDEBUGEVENT_indelay <= DBGC440UNCONDDEBUGEVENT_ipd after IN_DELAY;
	DCRPPCDMACK_indelay <= DCRPPCDMACK_ipd after IN_DELAY;
	DCRPPCDMDBUSIN_indelay <= DCRPPCDMDBUSIN_ipd after IN_DELAY;
	DCRPPCDMTIMEOUTWAIT_indelay <= DCRPPCDMTIMEOUTWAIT_ipd after IN_DELAY;
	DCRPPCDSABUS_indelay <= DCRPPCDSABUS_ipd after IN_DELAY;
	DCRPPCDSDBUSOUT_indelay <= DCRPPCDSDBUSOUT_ipd after IN_DELAY;
	DCRPPCDSREAD_indelay <= DCRPPCDSREAD_ipd after IN_DELAY;
	DCRPPCDSWRITE_indelay <= DCRPPCDSWRITE_ipd after IN_DELAY;
	EICC440CRITIRQ_indelay <= EICC440CRITIRQ_ipd after IN_DELAY;
	EICC440EXTIRQ_indelay <= EICC440EXTIRQ_ipd after IN_DELAY;
	FCMAPUCONFIRMINSTR_indelay <= FCMAPUCONFIRMINSTR_ipd after IN_DELAY;
	FCMAPUCR_indelay <= FCMAPUCR_ipd after IN_DELAY;
	FCMAPUDONE_indelay <= FCMAPUDONE_ipd after IN_DELAY;
	FCMAPUEXCEPTION_indelay <= FCMAPUEXCEPTION_ipd after IN_DELAY;
	FCMAPUFPSCRFEX_indelay <= FCMAPUFPSCRFEX_ipd after IN_DELAY;
	FCMAPURESULTVALID_indelay <= FCMAPURESULTVALID_ipd after IN_DELAY;
	FCMAPURESULT_indelay <= FCMAPURESULT_ipd after IN_DELAY;
	FCMAPUSLEEPNOTREADY_indelay <= FCMAPUSLEEPNOTREADY_ipd after IN_DELAY;
	FCMAPUSTOREDATA_indelay <= FCMAPUSTOREDATA_ipd after IN_DELAY;
	JTGC440TDI_indelay <= JTGC440TDI_ipd after IN_DELAY;
	JTGC440TMS_indelay <= JTGC440TMS_ipd after IN_DELAY;
	JTGC440TRSTNEG_indelay <= JTGC440TRSTNEG_ipd after IN_DELAY;
	LLDMA0RSTENGINEREQ_indelay <= LLDMA0RSTENGINEREQ_ipd after IN_DELAY;
	LLDMA0RXD_indelay <= LLDMA0RXD_ipd after IN_DELAY;
	LLDMA0RXEOFN_indelay <= LLDMA0RXEOFN_ipd after IN_DELAY;
	LLDMA0RXEOPN_indelay <= LLDMA0RXEOPN_ipd after IN_DELAY;
	LLDMA0RXREM_indelay <= LLDMA0RXREM_ipd after IN_DELAY;
	LLDMA0RXSOFN_indelay <= LLDMA0RXSOFN_ipd after IN_DELAY;
	LLDMA0RXSOPN_indelay <= LLDMA0RXSOPN_ipd after IN_DELAY;
	LLDMA0RXSRCRDYN_indelay <= LLDMA0RXSRCRDYN_ipd after IN_DELAY;
	LLDMA0TXDSTRDYN_indelay <= LLDMA0TXDSTRDYN_ipd after IN_DELAY;
	LLDMA1RSTENGINEREQ_indelay <= LLDMA1RSTENGINEREQ_ipd after IN_DELAY;
	LLDMA1RXD_indelay <= LLDMA1RXD_ipd after IN_DELAY;
	LLDMA1RXEOFN_indelay <= LLDMA1RXEOFN_ipd after IN_DELAY;
	LLDMA1RXEOPN_indelay <= LLDMA1RXEOPN_ipd after IN_DELAY;
	LLDMA1RXREM_indelay <= LLDMA1RXREM_ipd after IN_DELAY;
	LLDMA1RXSOFN_indelay <= LLDMA1RXSOFN_ipd after IN_DELAY;
	LLDMA1RXSOPN_indelay <= LLDMA1RXSOPN_ipd after IN_DELAY;
	LLDMA1RXSRCRDYN_indelay <= LLDMA1RXSRCRDYN_ipd after IN_DELAY;
	LLDMA1TXDSTRDYN_indelay <= LLDMA1TXDSTRDYN_ipd after IN_DELAY;
	LLDMA2RSTENGINEREQ_indelay <= LLDMA2RSTENGINEREQ_ipd after IN_DELAY;
	LLDMA2RXD_indelay <= LLDMA2RXD_ipd after IN_DELAY;
	LLDMA2RXEOFN_indelay <= LLDMA2RXEOFN_ipd after IN_DELAY;
	LLDMA2RXEOPN_indelay <= LLDMA2RXEOPN_ipd after IN_DELAY;
	LLDMA2RXREM_indelay <= LLDMA2RXREM_ipd after IN_DELAY;
	LLDMA2RXSOFN_indelay <= LLDMA2RXSOFN_ipd after IN_DELAY;
	LLDMA2RXSOPN_indelay <= LLDMA2RXSOPN_ipd after IN_DELAY;
	LLDMA2RXSRCRDYN_indelay <= LLDMA2RXSRCRDYN_ipd after IN_DELAY;
	LLDMA2TXDSTRDYN_indelay <= LLDMA2TXDSTRDYN_ipd after IN_DELAY;
	LLDMA3RSTENGINEREQ_indelay <= LLDMA3RSTENGINEREQ_ipd after IN_DELAY;
	LLDMA3RXD_indelay <= LLDMA3RXD_ipd after IN_DELAY;
	LLDMA3RXEOFN_indelay <= LLDMA3RXEOFN_ipd after IN_DELAY;
	LLDMA3RXEOPN_indelay <= LLDMA3RXEOPN_ipd after IN_DELAY;
	LLDMA3RXREM_indelay <= LLDMA3RXREM_ipd after IN_DELAY;
	LLDMA3RXSOFN_indelay <= LLDMA3RXSOFN_ipd after IN_DELAY;
	LLDMA3RXSOPN_indelay <= LLDMA3RXSOPN_ipd after IN_DELAY;
	LLDMA3RXSRCRDYN_indelay <= LLDMA3RXSRCRDYN_ipd after IN_DELAY;
	LLDMA3TXDSTRDYN_indelay <= LLDMA3TXDSTRDYN_ipd after IN_DELAY;
	MCMIADDRREADYTOACCEPT_indelay <= MCMIADDRREADYTOACCEPT_ipd after IN_DELAY;
	MCMIREADDATAERR_indelay <= MCMIREADDATAERR_ipd after IN_DELAY;
	MCMIREADDATAVALID_indelay <= MCMIREADDATAVALID_ipd after IN_DELAY;
	MCMIREADDATA_indelay <= MCMIREADDATA_ipd after IN_DELAY;
	PLBPPCMADDRACK_indelay <= PLBPPCMADDRACK_ipd after IN_DELAY;
	PLBPPCMMBUSY_indelay <= PLBPPCMMBUSY_ipd after IN_DELAY;
	PLBPPCMMIRQ_indelay <= PLBPPCMMIRQ_ipd after IN_DELAY;
	PLBPPCMMRDERR_indelay <= PLBPPCMMRDERR_ipd after IN_DELAY;
	PLBPPCMMWRERR_indelay <= PLBPPCMMWRERR_ipd after IN_DELAY;
	PLBPPCMRDBTERM_indelay <= PLBPPCMRDBTERM_ipd after IN_DELAY;
	PLBPPCMRDDACK_indelay <= PLBPPCMRDDACK_ipd after IN_DELAY;
	PLBPPCMRDDBUS_indelay <= PLBPPCMRDDBUS_ipd after IN_DELAY;
	PLBPPCMRDPENDPRI_indelay <= PLBPPCMRDPENDPRI_ipd after IN_DELAY;
	PLBPPCMRDPENDREQ_indelay <= PLBPPCMRDPENDREQ_ipd after IN_DELAY;
	PLBPPCMRDWDADDR_indelay <= PLBPPCMRDWDADDR_ipd after IN_DELAY;
	PLBPPCMREARBITRATE_indelay <= PLBPPCMREARBITRATE_ipd after IN_DELAY;
	PLBPPCMREQPRI_indelay <= PLBPPCMREQPRI_ipd after IN_DELAY;
	PLBPPCMSSIZE_indelay <= PLBPPCMSSIZE_ipd after IN_DELAY;
	PLBPPCMTIMEOUT_indelay <= PLBPPCMTIMEOUT_ipd after IN_DELAY;
	PLBPPCMWRBTERM_indelay <= PLBPPCMWRBTERM_ipd after IN_DELAY;
	PLBPPCMWRDACK_indelay <= PLBPPCMWRDACK_ipd after IN_DELAY;
	PLBPPCMWRPENDPRI_indelay <= PLBPPCMWRPENDPRI_ipd after IN_DELAY;
	PLBPPCMWRPENDREQ_indelay <= PLBPPCMWRPENDREQ_ipd after IN_DELAY;
	PLBPPCS0ABORT_indelay <= PLBPPCS0ABORT_ipd after IN_DELAY;
	PLBPPCS0ABUS_indelay <= PLBPPCS0ABUS_ipd after IN_DELAY;
	PLBPPCS0BE_indelay <= PLBPPCS0BE_ipd after IN_DELAY;
	PLBPPCS0BUSLOCK_indelay <= PLBPPCS0BUSLOCK_ipd after IN_DELAY;
	PLBPPCS0LOCKERR_indelay <= PLBPPCS0LOCKERR_ipd after IN_DELAY;
	PLBPPCS0MASTERID_indelay <= PLBPPCS0MASTERID_ipd after IN_DELAY;
	PLBPPCS0MSIZE_indelay <= PLBPPCS0MSIZE_ipd after IN_DELAY;
	PLBPPCS0PAVALID_indelay <= PLBPPCS0PAVALID_ipd after IN_DELAY;
	PLBPPCS0RDBURST_indelay <= PLBPPCS0RDBURST_ipd after IN_DELAY;
	PLBPPCS0RDPENDPRI_indelay <= PLBPPCS0RDPENDPRI_ipd after IN_DELAY;
	PLBPPCS0RDPENDREQ_indelay <= PLBPPCS0RDPENDREQ_ipd after IN_DELAY;
	PLBPPCS0RDPRIM_indelay <= PLBPPCS0RDPRIM_ipd after IN_DELAY;
	PLBPPCS0REQPRI_indelay <= PLBPPCS0REQPRI_ipd after IN_DELAY;
	PLBPPCS0RNW_indelay <= PLBPPCS0RNW_ipd after IN_DELAY;
	PLBPPCS0SAVALID_indelay <= PLBPPCS0SAVALID_ipd after IN_DELAY;
	PLBPPCS0SIZE_indelay <= PLBPPCS0SIZE_ipd after IN_DELAY;
	PLBPPCS0TATTRIBUTE_indelay <= PLBPPCS0TATTRIBUTE_ipd after IN_DELAY;
	PLBPPCS0TYPE_indelay <= PLBPPCS0TYPE_ipd after IN_DELAY;
	PLBPPCS0UABUS_indelay <= PLBPPCS0UABUS_ipd after IN_DELAY;
	PLBPPCS0WRBURST_indelay <= PLBPPCS0WRBURST_ipd after IN_DELAY;
	PLBPPCS0WRDBUS_indelay <= PLBPPCS0WRDBUS_ipd after IN_DELAY;
	PLBPPCS0WRPENDPRI_indelay <= PLBPPCS0WRPENDPRI_ipd after IN_DELAY;
	PLBPPCS0WRPENDREQ_indelay <= PLBPPCS0WRPENDREQ_ipd after IN_DELAY;
	PLBPPCS0WRPRIM_indelay <= PLBPPCS0WRPRIM_ipd after IN_DELAY;
	PLBPPCS1ABORT_indelay <= PLBPPCS1ABORT_ipd after IN_DELAY;
	PLBPPCS1ABUS_indelay <= PLBPPCS1ABUS_ipd after IN_DELAY;
	PLBPPCS1BE_indelay <= PLBPPCS1BE_ipd after IN_DELAY;
	PLBPPCS1BUSLOCK_indelay <= PLBPPCS1BUSLOCK_ipd after IN_DELAY;
	PLBPPCS1LOCKERR_indelay <= PLBPPCS1LOCKERR_ipd after IN_DELAY;
	PLBPPCS1MASTERID_indelay <= PLBPPCS1MASTERID_ipd after IN_DELAY;
	PLBPPCS1MSIZE_indelay <= PLBPPCS1MSIZE_ipd after IN_DELAY;
	PLBPPCS1PAVALID_indelay <= PLBPPCS1PAVALID_ipd after IN_DELAY;
	PLBPPCS1RDBURST_indelay <= PLBPPCS1RDBURST_ipd after IN_DELAY;
	PLBPPCS1RDPENDPRI_indelay <= PLBPPCS1RDPENDPRI_ipd after IN_DELAY;
	PLBPPCS1RDPENDREQ_indelay <= PLBPPCS1RDPENDREQ_ipd after IN_DELAY;
	PLBPPCS1RDPRIM_indelay <= PLBPPCS1RDPRIM_ipd after IN_DELAY;
	PLBPPCS1REQPRI_indelay <= PLBPPCS1REQPRI_ipd after IN_DELAY;
	PLBPPCS1RNW_indelay <= PLBPPCS1RNW_ipd after IN_DELAY;
	PLBPPCS1SAVALID_indelay <= PLBPPCS1SAVALID_ipd after IN_DELAY;
	PLBPPCS1SIZE_indelay <= PLBPPCS1SIZE_ipd after IN_DELAY;
	PLBPPCS1TATTRIBUTE_indelay <= PLBPPCS1TATTRIBUTE_ipd after IN_DELAY;
	PLBPPCS1TYPE_indelay <= PLBPPCS1TYPE_ipd after IN_DELAY;
	PLBPPCS1UABUS_indelay <= PLBPPCS1UABUS_ipd after IN_DELAY;
	PLBPPCS1WRBURST_indelay <= PLBPPCS1WRBURST_ipd after IN_DELAY;
	PLBPPCS1WRDBUS_indelay <= PLBPPCS1WRDBUS_ipd after IN_DELAY;
	PLBPPCS1WRPENDPRI_indelay <= PLBPPCS1WRPENDPRI_ipd after IN_DELAY;
	PLBPPCS1WRPENDREQ_indelay <= PLBPPCS1WRPENDREQ_ipd after IN_DELAY;
	PLBPPCS1WRPRIM_indelay <= PLBPPCS1WRPRIM_ipd after IN_DELAY;
	RSTC440RESETCHIP_indelay <= RSTC440RESETCHIP_ipd after IN_DELAY;
	RSTC440RESETCORE_indelay <= RSTC440RESETCORE_ipd after IN_DELAY;
	RSTC440RESETSYSTEM_indelay <= RSTC440RESETSYSTEM_ipd after IN_DELAY;
	TIEC440DCURDLDCACHEPLBPRIO_indelay <= TIEC440DCURDLDCACHEPLBPRIO_ipd after IN_DELAY;
	TIEC440DCURDNONCACHEPLBPRIO_indelay <= TIEC440DCURDNONCACHEPLBPRIO_ipd after IN_DELAY;
	TIEC440DCURDTOUCHPLBPRIO_indelay <= TIEC440DCURDTOUCHPLBPRIO_ipd after IN_DELAY;
	TIEC440DCURDURGENTPLBPRIO_indelay <= TIEC440DCURDURGENTPLBPRIO_ipd after IN_DELAY;
	TIEC440DCUWRFLUSHPLBPRIO_indelay <= TIEC440DCUWRFLUSHPLBPRIO_ipd after IN_DELAY;
	TIEC440DCUWRSTOREPLBPRIO_indelay <= TIEC440DCUWRSTOREPLBPRIO_ipd after IN_DELAY;
	TIEC440DCUWRURGENTPLBPRIO_indelay <= TIEC440DCUWRURGENTPLBPRIO_ipd after IN_DELAY;
	TIEC440ENDIANRESET_indelay <= TIEC440ENDIANRESET_ipd after IN_DELAY;
	TIEC440ERPNRESET_indelay <= TIEC440ERPNRESET_ipd after IN_DELAY;
	TIEC440ICURDFETCHPLBPRIO_indelay <= TIEC440ICURDFETCHPLBPRIO_ipd after IN_DELAY;
	TIEC440ICURDSPECPLBPRIO_indelay <= TIEC440ICURDSPECPLBPRIO_ipd after IN_DELAY;
	TIEC440ICURDTOUCHPLBPRIO_indelay <= TIEC440ICURDTOUCHPLBPRIO_ipd after IN_DELAY;
	TIEC440PIR_indelay <= TIEC440PIR_ipd after IN_DELAY;
	TIEC440PVR_indelay <= TIEC440PVR_ipd after IN_DELAY;
	TIEC440USERRESET_indelay <= TIEC440USERRESET_ipd after IN_DELAY;
	TIEDCRBASEADDR_indelay <= TIEDCRBASEADDR_ipd after IN_DELAY;
	TRCC440TRACEDISABLE_indelay <= TRCC440TRACEDISABLE_ipd after IN_DELAY;
	TRCC440TRIGGEREVENTIN_indelay <= TRCC440TRIGGEREVENTIN_ipd after IN_DELAY;


	ppc440_swift_1 : PPC440_SWIFT
	port map (
	APU_CONTROL  =>  APU_CONTROL_BINARY,
	APU_UDI0  =>  APU_UDI0_BINARY,
	APU_UDI1  =>  APU_UDI1_BINARY,
	APU_UDI10  =>  APU_UDI10_BINARY,
	APU_UDI11  =>  APU_UDI11_BINARY,
	APU_UDI12  =>  APU_UDI12_BINARY,
	APU_UDI13  =>  APU_UDI13_BINARY,
	APU_UDI14  =>  APU_UDI14_BINARY,
	APU_UDI15  =>  APU_UDI15_BINARY,
	APU_UDI2  =>  APU_UDI2_BINARY,
	APU_UDI3  =>  APU_UDI3_BINARY,
	APU_UDI4  =>  APU_UDI4_BINARY,
	APU_UDI5  =>  APU_UDI5_BINARY,
	APU_UDI6  =>  APU_UDI6_BINARY,
	APU_UDI7  =>  APU_UDI7_BINARY,
	APU_UDI8  =>  APU_UDI8_BINARY,
	APU_UDI9  =>  APU_UDI9_BINARY,
	CLOCK_DELAY  =>  CLOCK_DELAY_BINARY,
	DCR_AUTOLOCK_ENABLE  =>  DCR_AUTOLOCK_ENABLE_BINARY,
	DMA0_CONTROL  =>  DMA0_CONTROL_BINARY,
	DMA0_RXCHANNELCTRL  =>  DMA0_RXCHANNELCTRL_BINARY,
	DMA0_RXIRQTIMER  =>  DMA0_RXIRQTIMER_BINARY,
	DMA0_TXCHANNELCTRL  =>  DMA0_TXCHANNELCTRL_BINARY,
	DMA0_TXIRQTIMER  =>  DMA0_TXIRQTIMER_BINARY,
	DMA1_CONTROL  =>  DMA1_CONTROL_BINARY,
	DMA1_RXCHANNELCTRL  =>  DMA1_RXCHANNELCTRL_BINARY,
	DMA1_RXIRQTIMER  =>  DMA1_RXIRQTIMER_BINARY,
	DMA1_TXCHANNELCTRL  =>  DMA1_TXCHANNELCTRL_BINARY,
	DMA1_TXIRQTIMER  =>  DMA1_TXIRQTIMER_BINARY,
	DMA2_CONTROL  =>  DMA2_CONTROL_BINARY,
	DMA2_RXCHANNELCTRL  =>  DMA2_RXCHANNELCTRL_BINARY,
	DMA2_RXIRQTIMER  =>  DMA2_RXIRQTIMER_BINARY,
	DMA2_TXCHANNELCTRL  =>  DMA2_TXCHANNELCTRL_BINARY,
	DMA2_TXIRQTIMER  =>  DMA2_TXIRQTIMER_BINARY,
	DMA3_CONTROL  =>  DMA3_CONTROL_BINARY,
	DMA3_RXCHANNELCTRL  =>  DMA3_RXCHANNELCTRL_BINARY,
	DMA3_RXIRQTIMER  =>  DMA3_RXIRQTIMER_BINARY,
	DMA3_TXCHANNELCTRL  =>  DMA3_TXCHANNELCTRL_BINARY,
	DMA3_TXIRQTIMER  =>  DMA3_TXIRQTIMER_BINARY,
	INTERCONNECT_IMASK  =>  INTERCONNECT_IMASK_BINARY,
	INTERCONNECT_TMPL_SEL  =>  INTERCONNECT_TMPL_SEL_BINARY,
	MI_ARBCONFIG  =>  MI_ARBCONFIG_BINARY,
	MI_BANKCONFLICT_MASK  =>  MI_BANKCONFLICT_MASK_BINARY,
	MI_CONTROL  =>  MI_CONTROL_BINARY,
	MI_ROWCONFLICT_MASK  =>  MI_ROWCONFLICT_MASK_BINARY,
	PPCDM_ASYNCMODE  =>  PPCDM_ASYNCMODE_BINARY,
	PPCDS_ASYNCMODE  =>  PPCDS_ASYNCMODE_BINARY,
	PPCM_ARBCONFIG  =>  PPCM_ARBCONFIG_BINARY,
	PPCM_CONTROL  =>  PPCM_CONTROL_BINARY,
	PPCM_COUNTER  =>  PPCM_COUNTER_BINARY,
	PPCS0_ADDRMAP_TMPL0  =>  PPCS0_ADDRMAP_TMPL0_BINARY,
	PPCS0_ADDRMAP_TMPL1  =>  PPCS0_ADDRMAP_TMPL1_BINARY,
	PPCS0_ADDRMAP_TMPL2  =>  PPCS0_ADDRMAP_TMPL2_BINARY,
	PPCS0_ADDRMAP_TMPL3  =>  PPCS0_ADDRMAP_TMPL3_BINARY,
	PPCS0_CONTROL  =>  PPCS0_CONTROL_BINARY,
	PPCS0_WIDTH_128N64  =>  PPCS0_WIDTH_128N64_BINARY,
	PPCS1_ADDRMAP_TMPL0  =>  PPCS1_ADDRMAP_TMPL0_BINARY,
	PPCS1_ADDRMAP_TMPL1  =>  PPCS1_ADDRMAP_TMPL1_BINARY,
	PPCS1_ADDRMAP_TMPL2  =>  PPCS1_ADDRMAP_TMPL2_BINARY,
	PPCS1_ADDRMAP_TMPL3  =>  PPCS1_ADDRMAP_TMPL3_BINARY,
	PPCS1_CONTROL  =>  PPCS1_CONTROL_BINARY,
	PPCS1_WIDTH_128N64  =>  PPCS1_WIDTH_128N64_BINARY,
	XBAR_ADDRMAP_TMPL0  =>  XBAR_ADDRMAP_TMPL0_BINARY,
	XBAR_ADDRMAP_TMPL1  =>  XBAR_ADDRMAP_TMPL1_BINARY,
	XBAR_ADDRMAP_TMPL2  =>  XBAR_ADDRMAP_TMPL2_BINARY,
	XBAR_ADDRMAP_TMPL3  =>  XBAR_ADDRMAP_TMPL3_BINARY,

	APUFCMDECFPUOP  =>  APUFCMDECFPUOP_outdelay,
	APUFCMDECLDSTXFERSIZE  =>  APUFCMDECLDSTXFERSIZE_outdelay,
	APUFCMDECLOAD  =>  APUFCMDECLOAD_outdelay,
	APUFCMDECNONAUTON  =>  APUFCMDECNONAUTON_outdelay,
	APUFCMDECSTORE  =>  APUFCMDECSTORE_outdelay,
	APUFCMDECUDI  =>  APUFCMDECUDI_outdelay,
	APUFCMDECUDIVALID  =>  APUFCMDECUDIVALID_outdelay,
	APUFCMENDIAN  =>  APUFCMENDIAN_outdelay,
	APUFCMFLUSH  =>  APUFCMFLUSH_outdelay,
	APUFCMINSTRUCTION  =>  APUFCMINSTRUCTION_outdelay,
	APUFCMINSTRVALID  =>  APUFCMINSTRVALID_outdelay,
	APUFCMLOADBYTEADDR  =>  APUFCMLOADBYTEADDR_outdelay,
	APUFCMLOADDATA  =>  APUFCMLOADDATA_outdelay,
	APUFCMLOADDVALID  =>  APUFCMLOADDVALID_outdelay,
	APUFCMMSRFE0  =>  APUFCMMSRFE0_outdelay,
	APUFCMMSRFE1  =>  APUFCMMSRFE1_outdelay,
	APUFCMNEXTINSTRREADY  =>  APUFCMNEXTINSTRREADY_outdelay,
	APUFCMOPERANDVALID  =>  APUFCMOPERANDVALID_outdelay,
	APUFCMRADATA  =>  APUFCMRADATA_outdelay,
	APUFCMRBDATA  =>  APUFCMRBDATA_outdelay,
	APUFCMWRITEBACKOK  =>  APUFCMWRITEBACKOK_outdelay,
	C440CPMCORESLEEPREQ  =>  C440CPMCORESLEEPREQ_outdelay,
	C440CPMDECIRPTREQ  =>  C440CPMDECIRPTREQ_outdelay,
	C440CPMFITIRPTREQ  =>  C440CPMFITIRPTREQ_outdelay,
	C440CPMMSRCE  =>  C440CPMMSRCE_outdelay,
	C440CPMMSREE  =>  C440CPMMSREE_outdelay,
	C440CPMTIMERRESETREQ  =>  C440CPMTIMERRESETREQ_outdelay,
	C440CPMWDIRPTREQ  =>  C440CPMWDIRPTREQ_outdelay,
	C440DBGSYSTEMCONTROL  =>  C440DBGSYSTEMCONTROL_outdelay,
	C440JTGTDO  =>  C440JTGTDO_outdelay,
	C440JTGTDOEN  =>  C440JTGTDOEN_outdelay,
	C440MACHINECHECK  =>  C440MACHINECHECK_outdelay,
	C440RSTCHIPRESETREQ  =>  C440RSTCHIPRESETREQ_outdelay,
	C440RSTCORERESETREQ  =>  C440RSTCORERESETREQ_outdelay,
	C440RSTSYSTEMRESETREQ  =>  C440RSTSYSTEMRESETREQ_outdelay,
	C440TRCBRANCHSTATUS  =>  C440TRCBRANCHSTATUS_outdelay,
	C440TRCCYCLE  =>  C440TRCCYCLE_outdelay,
	C440TRCEXECUTIONSTATUS  =>  C440TRCEXECUTIONSTATUS_outdelay,
	C440TRCTRACESTATUS  =>  C440TRCTRACESTATUS_outdelay,
	C440TRCTRIGGEREVENTOUT  =>  C440TRCTRIGGEREVENTOUT_outdelay,
	C440TRCTRIGGEREVENTTYPE  =>  C440TRCTRIGGEREVENTTYPE_outdelay,
	DMA0LLRSTENGINEACK  =>  DMA0LLRSTENGINEACK_outdelay,
	DMA0LLRXDSTRDYN  =>  DMA0LLRXDSTRDYN_outdelay,
	DMA0LLTXD  =>  DMA0LLTXD_outdelay,
	DMA0LLTXEOFN  =>  DMA0LLTXEOFN_outdelay,
	DMA0LLTXEOPN  =>  DMA0LLTXEOPN_outdelay,
	DMA0LLTXREM  =>  DMA0LLTXREM_outdelay,
	DMA0LLTXSOFN  =>  DMA0LLTXSOFN_outdelay,
	DMA0LLTXSOPN  =>  DMA0LLTXSOPN_outdelay,
	DMA0LLTXSRCRDYN  =>  DMA0LLTXSRCRDYN_outdelay,
	DMA0RXIRQ  =>  DMA0RXIRQ_outdelay,
	DMA0TXIRQ  =>  DMA0TXIRQ_outdelay,
	DMA1LLRSTENGINEACK  =>  DMA1LLRSTENGINEACK_outdelay,
	DMA1LLRXDSTRDYN  =>  DMA1LLRXDSTRDYN_outdelay,
	DMA1LLTXD  =>  DMA1LLTXD_outdelay,
	DMA1LLTXEOFN  =>  DMA1LLTXEOFN_outdelay,
	DMA1LLTXEOPN  =>  DMA1LLTXEOPN_outdelay,
	DMA1LLTXREM  =>  DMA1LLTXREM_outdelay,
	DMA1LLTXSOFN  =>  DMA1LLTXSOFN_outdelay,
	DMA1LLTXSOPN  =>  DMA1LLTXSOPN_outdelay,
	DMA1LLTXSRCRDYN  =>  DMA1LLTXSRCRDYN_outdelay,
	DMA1RXIRQ  =>  DMA1RXIRQ_outdelay,
	DMA1TXIRQ  =>  DMA1TXIRQ_outdelay,
	DMA2LLRSTENGINEACK  =>  DMA2LLRSTENGINEACK_outdelay,
	DMA2LLRXDSTRDYN  =>  DMA2LLRXDSTRDYN_outdelay,
	DMA2LLTXD  =>  DMA2LLTXD_outdelay,
	DMA2LLTXEOFN  =>  DMA2LLTXEOFN_outdelay,
	DMA2LLTXEOPN  =>  DMA2LLTXEOPN_outdelay,
	DMA2LLTXREM  =>  DMA2LLTXREM_outdelay,
	DMA2LLTXSOFN  =>  DMA2LLTXSOFN_outdelay,
	DMA2LLTXSOPN  =>  DMA2LLTXSOPN_outdelay,
	DMA2LLTXSRCRDYN  =>  DMA2LLTXSRCRDYN_outdelay,
	DMA2RXIRQ  =>  DMA2RXIRQ_outdelay,
	DMA2TXIRQ  =>  DMA2TXIRQ_outdelay,
	DMA3LLRSTENGINEACK  =>  DMA3LLRSTENGINEACK_outdelay,
	DMA3LLRXDSTRDYN  =>  DMA3LLRXDSTRDYN_outdelay,
	DMA3LLTXD  =>  DMA3LLTXD_outdelay,
	DMA3LLTXEOFN  =>  DMA3LLTXEOFN_outdelay,
	DMA3LLTXEOPN  =>  DMA3LLTXEOPN_outdelay,
	DMA3LLTXREM  =>  DMA3LLTXREM_outdelay,
	DMA3LLTXSOFN  =>  DMA3LLTXSOFN_outdelay,
	DMA3LLTXSOPN  =>  DMA3LLTXSOPN_outdelay,
	DMA3LLTXSRCRDYN  =>  DMA3LLTXSRCRDYN_outdelay,
	DMA3RXIRQ  =>  DMA3RXIRQ_outdelay,
	DMA3TXIRQ  =>  DMA3TXIRQ_outdelay,
	MIMCADDRESS  =>  MIMCADDRESS_outdelay,
	MIMCADDRESSVALID  =>  MIMCADDRESSVALID_outdelay,
	MIMCBANKCONFLICT  =>  MIMCBANKCONFLICT_outdelay,
	MIMCBYTEENABLE  =>  MIMCBYTEENABLE_outdelay,
	MIMCREADNOTWRITE  =>  MIMCREADNOTWRITE_outdelay,
	MIMCROWCONFLICT  =>  MIMCROWCONFLICT_outdelay,
	MIMCWRITEDATA  =>  MIMCWRITEDATA_outdelay,
	MIMCWRITEDATAVALID  =>  MIMCWRITEDATAVALID_outdelay,
	PPCCPMINTERCONNECTBUSY  =>  PPCCPMINTERCONNECTBUSY_outdelay,
	PPCDMDCRABUS  =>  PPCDMDCRABUS_outdelay,
	PPCDMDCRDBUSOUT  =>  PPCDMDCRDBUSOUT_outdelay,
	PPCDMDCRREAD  =>  PPCDMDCRREAD_outdelay,
	PPCDMDCRUABUS  =>  PPCDMDCRUABUS_outdelay,
	PPCDMDCRWRITE  =>  PPCDMDCRWRITE_outdelay,
	PPCDSDCRACK  =>  PPCDSDCRACK_outdelay,
	PPCDSDCRDBUSIN  =>  PPCDSDCRDBUSIN_outdelay,
	PPCDSDCRTIMEOUTWAIT  =>  PPCDSDCRTIMEOUTWAIT_outdelay,
	PPCEICINTERCONNECTIRQ  =>  PPCEICINTERCONNECTIRQ_outdelay,
	PPCMPLBABORT  =>  PPCMPLBABORT_outdelay,
	PPCMPLBABUS  =>  PPCMPLBABUS_outdelay,
	PPCMPLBBE  =>  PPCMPLBBE_outdelay,
	PPCMPLBBUSLOCK  =>  PPCMPLBBUSLOCK_outdelay,
	PPCMPLBLOCKERR  =>  PPCMPLBLOCKERR_outdelay,
	PPCMPLBPRIORITY  =>  PPCMPLBPRIORITY_outdelay,
	PPCMPLBRDBURST  =>  PPCMPLBRDBURST_outdelay,
	PPCMPLBREQUEST  =>  PPCMPLBREQUEST_outdelay,
	PPCMPLBRNW  =>  PPCMPLBRNW_outdelay,
	PPCMPLBSIZE  =>  PPCMPLBSIZE_outdelay,
	PPCMPLBTATTRIBUTE  =>  PPCMPLBTATTRIBUTE_outdelay,
	PPCMPLBTYPE  =>  PPCMPLBTYPE_outdelay,
	PPCMPLBUABUS  =>  PPCMPLBUABUS_outdelay,
	PPCMPLBWRBURST  =>  PPCMPLBWRBURST_outdelay,
	PPCMPLBWRDBUS  =>  PPCMPLBWRDBUS_outdelay,
	PPCS0PLBADDRACK  =>  PPCS0PLBADDRACK_outdelay,
	PPCS0PLBMBUSY  =>  PPCS0PLBMBUSY_outdelay,
	PPCS0PLBMIRQ  =>  PPCS0PLBMIRQ_outdelay,
	PPCS0PLBMRDERR  =>  PPCS0PLBMRDERR_outdelay,
	PPCS0PLBMWRERR  =>  PPCS0PLBMWRERR_outdelay,
	PPCS0PLBRDBTERM  =>  PPCS0PLBRDBTERM_outdelay,
	PPCS0PLBRDCOMP  =>  PPCS0PLBRDCOMP_outdelay,
	PPCS0PLBRDDACK  =>  PPCS0PLBRDDACK_outdelay,
	PPCS0PLBRDDBUS  =>  PPCS0PLBRDDBUS_outdelay,
	PPCS0PLBRDWDADDR  =>  PPCS0PLBRDWDADDR_outdelay,
	PPCS0PLBREARBITRATE  =>  PPCS0PLBREARBITRATE_outdelay,
	PPCS0PLBSSIZE  =>  PPCS0PLBSSIZE_outdelay,
	PPCS0PLBWAIT  =>  PPCS0PLBWAIT_outdelay,
	PPCS0PLBWRBTERM  =>  PPCS0PLBWRBTERM_outdelay,
	PPCS0PLBWRCOMP  =>  PPCS0PLBWRCOMP_outdelay,
	PPCS0PLBWRDACK  =>  PPCS0PLBWRDACK_outdelay,
	PPCS1PLBADDRACK  =>  PPCS1PLBADDRACK_outdelay,
	PPCS1PLBMBUSY  =>  PPCS1PLBMBUSY_outdelay,
	PPCS1PLBMIRQ  =>  PPCS1PLBMIRQ_outdelay,
	PPCS1PLBMRDERR  =>  PPCS1PLBMRDERR_outdelay,
	PPCS1PLBMWRERR  =>  PPCS1PLBMWRERR_outdelay,
	PPCS1PLBRDBTERM  =>  PPCS1PLBRDBTERM_outdelay,
	PPCS1PLBRDCOMP  =>  PPCS1PLBRDCOMP_outdelay,
	PPCS1PLBRDDACK  =>  PPCS1PLBRDDACK_outdelay,
	PPCS1PLBRDDBUS  =>  PPCS1PLBRDDBUS_outdelay,
	PPCS1PLBRDWDADDR  =>  PPCS1PLBRDWDADDR_outdelay,
	PPCS1PLBREARBITRATE  =>  PPCS1PLBREARBITRATE_outdelay,
	PPCS1PLBSSIZE  =>  PPCS1PLBSSIZE_outdelay,
	PPCS1PLBWAIT  =>  PPCS1PLBWAIT_outdelay,
	PPCS1PLBWRBTERM  =>  PPCS1PLBWRBTERM_outdelay,
	PPCS1PLBWRCOMP  =>  PPCS1PLBWRCOMP_outdelay,
	PPCS1PLBWRDACK  =>  PPCS1PLBWRDACK_outdelay,

	CPMC440CLK  =>  CPMC440CLK_indelay,
	CPMC440CLKEN  =>  CPMC440CLKEN_indelay,
	CPMC440CORECLOCKINACTIVE  =>  CPMC440CORECLOCKINACTIVE_indelay,
	CPMC440TIMERCLOCK  =>  CPMC440TIMERCLOCK_indelay,
	CPMDCRCLK  =>  CPMDCRCLK_indelay,
	CPMDMA0LLCLK  =>  CPMDMA0LLCLK_indelay,
	CPMDMA1LLCLK  =>  CPMDMA1LLCLK_indelay,
	CPMDMA2LLCLK  =>  CPMDMA2LLCLK_indelay,
	CPMDMA3LLCLK  =>  CPMDMA3LLCLK_indelay,
	CPMFCMCLK  =>  CPMFCMCLK_indelay,
	CPMINTERCONNECTCLK  =>  CPMINTERCONNECTCLK_indelay,
	CPMINTERCONNECTCLKEN  =>  CPMINTERCONNECTCLKEN_indelay,
	CPMINTERCONNECTCLKNTO1  =>  CPMINTERCONNECTCLKNTO1_indelay,
	CPMMCCLK  =>  CPMMCCLK_indelay,
	CPMPPCMPLBCLK  =>  CPMPPCMPLBCLK_indelay,
	CPMPPCS0PLBCLK  =>  CPMPPCS0PLBCLK_indelay,
	CPMPPCS1PLBCLK  =>  CPMPPCS1PLBCLK_indelay,
	DBGC440DEBUGHALT  =>  DBGC440DEBUGHALT_indelay,
	DBGC440SYSTEMSTATUS  =>  DBGC440SYSTEMSTATUS_indelay,
	DBGC440UNCONDDEBUGEVENT  =>  DBGC440UNCONDDEBUGEVENT_indelay,
	DCRPPCDMACK  =>  DCRPPCDMACK_indelay,
	DCRPPCDMDBUSIN  =>  DCRPPCDMDBUSIN_indelay,
	DCRPPCDMTIMEOUTWAIT  =>  DCRPPCDMTIMEOUTWAIT_indelay,
	DCRPPCDSABUS  =>  DCRPPCDSABUS_indelay,
	DCRPPCDSDBUSOUT  =>  DCRPPCDSDBUSOUT_indelay,
	DCRPPCDSREAD  =>  DCRPPCDSREAD_indelay,
	DCRPPCDSWRITE  =>  DCRPPCDSWRITE_indelay,
	EICC440CRITIRQ  =>  EICC440CRITIRQ_indelay,
	EICC440EXTIRQ  =>  EICC440EXTIRQ_indelay,
	FCMAPUCONFIRMINSTR  =>  FCMAPUCONFIRMINSTR_indelay,
	FCMAPUCR  =>  FCMAPUCR_indelay,
	FCMAPUDONE  =>  FCMAPUDONE_indelay,
	FCMAPUEXCEPTION  =>  FCMAPUEXCEPTION_indelay,
	FCMAPUFPSCRFEX  =>  FCMAPUFPSCRFEX_indelay,
	FCMAPURESULT  =>  FCMAPURESULT_indelay,
	FCMAPURESULTVALID  =>  FCMAPURESULTVALID_indelay,
	FCMAPUSLEEPNOTREADY  =>  FCMAPUSLEEPNOTREADY_indelay,
	FCMAPUSTOREDATA  =>  FCMAPUSTOREDATA_indelay,
	GSR  =>  GSR,
	JTGC440TCK  =>  JTGC440TCK_indelay,
	JTGC440TDI  =>  JTGC440TDI_indelay,
	JTGC440TMS  =>  JTGC440TMS_indelay,
	JTGC440TRSTNEG  =>  JTGC440TRSTNEG_indelay,
	LLDMA0RSTENGINEREQ  =>  LLDMA0RSTENGINEREQ_indelay,
	LLDMA0RXD  =>  LLDMA0RXD_indelay,
	LLDMA0RXEOFN  =>  LLDMA0RXEOFN_indelay,
	LLDMA0RXEOPN  =>  LLDMA0RXEOPN_indelay,
	LLDMA0RXREM  =>  LLDMA0RXREM_indelay,
	LLDMA0RXSOFN  =>  LLDMA0RXSOFN_indelay,
	LLDMA0RXSOPN  =>  LLDMA0RXSOPN_indelay,
	LLDMA0RXSRCRDYN  =>  LLDMA0RXSRCRDYN_indelay,
	LLDMA0TXDSTRDYN  =>  LLDMA0TXDSTRDYN_indelay,
	LLDMA1RSTENGINEREQ  =>  LLDMA1RSTENGINEREQ_indelay,
	LLDMA1RXD  =>  LLDMA1RXD_indelay,
	LLDMA1RXEOFN  =>  LLDMA1RXEOFN_indelay,
	LLDMA1RXEOPN  =>  LLDMA1RXEOPN_indelay,
	LLDMA1RXREM  =>  LLDMA1RXREM_indelay,
	LLDMA1RXSOFN  =>  LLDMA1RXSOFN_indelay,
	LLDMA1RXSOPN  =>  LLDMA1RXSOPN_indelay,
	LLDMA1RXSRCRDYN  =>  LLDMA1RXSRCRDYN_indelay,
	LLDMA1TXDSTRDYN  =>  LLDMA1TXDSTRDYN_indelay,
	LLDMA2RSTENGINEREQ  =>  LLDMA2RSTENGINEREQ_indelay,
	LLDMA2RXD  =>  LLDMA2RXD_indelay,
	LLDMA2RXEOFN  =>  LLDMA2RXEOFN_indelay,
	LLDMA2RXEOPN  =>  LLDMA2RXEOPN_indelay,
	LLDMA2RXREM  =>  LLDMA2RXREM_indelay,
	LLDMA2RXSOFN  =>  LLDMA2RXSOFN_indelay,
	LLDMA2RXSOPN  =>  LLDMA2RXSOPN_indelay,
	LLDMA2RXSRCRDYN  =>  LLDMA2RXSRCRDYN_indelay,
	LLDMA2TXDSTRDYN  =>  LLDMA2TXDSTRDYN_indelay,
	LLDMA3RSTENGINEREQ  =>  LLDMA3RSTENGINEREQ_indelay,
	LLDMA3RXD  =>  LLDMA3RXD_indelay,
	LLDMA3RXEOFN  =>  LLDMA3RXEOFN_indelay,
	LLDMA3RXEOPN  =>  LLDMA3RXEOPN_indelay,
	LLDMA3RXREM  =>  LLDMA3RXREM_indelay,
	LLDMA3RXSOFN  =>  LLDMA3RXSOFN_indelay,
	LLDMA3RXSOPN  =>  LLDMA3RXSOPN_indelay,
	LLDMA3RXSRCRDYN  =>  LLDMA3RXSRCRDYN_indelay,
	LLDMA3TXDSTRDYN  =>  LLDMA3TXDSTRDYN_indelay,
	MCMIADDRREADYTOACCEPT  =>  MCMIADDRREADYTOACCEPT_indelay,
	MCMIREADDATA  =>  MCMIREADDATA_indelay,
	MCMIREADDATAERR  =>  MCMIREADDATAERR_indelay,
	MCMIREADDATAVALID  =>  MCMIREADDATAVALID_indelay,
	PLBPPCMADDRACK  =>  PLBPPCMADDRACK_indelay,
	PLBPPCMMBUSY  =>  PLBPPCMMBUSY_indelay,
	PLBPPCMMIRQ  =>  PLBPPCMMIRQ_indelay,
	PLBPPCMMRDERR  =>  PLBPPCMMRDERR_indelay,
	PLBPPCMMWRERR  =>  PLBPPCMMWRERR_indelay,
	PLBPPCMRDBTERM  =>  PLBPPCMRDBTERM_indelay,
	PLBPPCMRDDACK  =>  PLBPPCMRDDACK_indelay,
	PLBPPCMRDDBUS  =>  PLBPPCMRDDBUS_indelay,
	PLBPPCMRDPENDPRI  =>  PLBPPCMRDPENDPRI_indelay,
	PLBPPCMRDPENDREQ  =>  PLBPPCMRDPENDREQ_indelay,
	PLBPPCMRDWDADDR  =>  PLBPPCMRDWDADDR_indelay,
	PLBPPCMREARBITRATE  =>  PLBPPCMREARBITRATE_indelay,
	PLBPPCMREQPRI  =>  PLBPPCMREQPRI_indelay,
	PLBPPCMSSIZE  =>  PLBPPCMSSIZE_indelay,
	PLBPPCMTIMEOUT  =>  PLBPPCMTIMEOUT_indelay,
	PLBPPCMWRBTERM  =>  PLBPPCMWRBTERM_indelay,
	PLBPPCMWRDACK  =>  PLBPPCMWRDACK_indelay,
	PLBPPCMWRPENDPRI  =>  PLBPPCMWRPENDPRI_indelay,
	PLBPPCMWRPENDREQ  =>  PLBPPCMWRPENDREQ_indelay,
	PLBPPCS0ABORT  =>  PLBPPCS0ABORT_indelay,
	PLBPPCS0ABUS  =>  PLBPPCS0ABUS_indelay,
	PLBPPCS0BE  =>  PLBPPCS0BE_indelay,
	PLBPPCS0BUSLOCK  =>  PLBPPCS0BUSLOCK_indelay,
	PLBPPCS0LOCKERR  =>  PLBPPCS0LOCKERR_indelay,
	PLBPPCS0MASTERID  =>  PLBPPCS0MASTERID_indelay,
	PLBPPCS0MSIZE  =>  PLBPPCS0MSIZE_indelay,
	PLBPPCS0PAVALID  =>  PLBPPCS0PAVALID_indelay,
	PLBPPCS0RDBURST  =>  PLBPPCS0RDBURST_indelay,
	PLBPPCS0RDPENDPRI  =>  PLBPPCS0RDPENDPRI_indelay,
	PLBPPCS0RDPENDREQ  =>  PLBPPCS0RDPENDREQ_indelay,
	PLBPPCS0RDPRIM  =>  PLBPPCS0RDPRIM_indelay,
	PLBPPCS0REQPRI  =>  PLBPPCS0REQPRI_indelay,
	PLBPPCS0RNW  =>  PLBPPCS0RNW_indelay,
	PLBPPCS0SAVALID  =>  PLBPPCS0SAVALID_indelay,
	PLBPPCS0SIZE  =>  PLBPPCS0SIZE_indelay,
	PLBPPCS0TATTRIBUTE  =>  PLBPPCS0TATTRIBUTE_indelay,
	PLBPPCS0TYPE  =>  PLBPPCS0TYPE_indelay,
	PLBPPCS0UABUS  =>  PLBPPCS0UABUS_indelay,
	PLBPPCS0WRBURST  =>  PLBPPCS0WRBURST_indelay,
	PLBPPCS0WRDBUS  =>  PLBPPCS0WRDBUS_indelay,
	PLBPPCS0WRPENDPRI  =>  PLBPPCS0WRPENDPRI_indelay,
	PLBPPCS0WRPENDREQ  =>  PLBPPCS0WRPENDREQ_indelay,
	PLBPPCS0WRPRIM  =>  PLBPPCS0WRPRIM_indelay,
	PLBPPCS1ABORT  =>  PLBPPCS1ABORT_indelay,
	PLBPPCS1ABUS  =>  PLBPPCS1ABUS_indelay,
	PLBPPCS1BE  =>  PLBPPCS1BE_indelay,
	PLBPPCS1BUSLOCK  =>  PLBPPCS1BUSLOCK_indelay,
	PLBPPCS1LOCKERR  =>  PLBPPCS1LOCKERR_indelay,
	PLBPPCS1MASTERID  =>  PLBPPCS1MASTERID_indelay,
	PLBPPCS1MSIZE  =>  PLBPPCS1MSIZE_indelay,
	PLBPPCS1PAVALID  =>  PLBPPCS1PAVALID_indelay,
	PLBPPCS1RDBURST  =>  PLBPPCS1RDBURST_indelay,
	PLBPPCS1RDPENDPRI  =>  PLBPPCS1RDPENDPRI_indelay,
	PLBPPCS1RDPENDREQ  =>  PLBPPCS1RDPENDREQ_indelay,
	PLBPPCS1RDPRIM  =>  PLBPPCS1RDPRIM_indelay,
	PLBPPCS1REQPRI  =>  PLBPPCS1REQPRI_indelay,
	PLBPPCS1RNW  =>  PLBPPCS1RNW_indelay,
	PLBPPCS1SAVALID  =>  PLBPPCS1SAVALID_indelay,
	PLBPPCS1SIZE  =>  PLBPPCS1SIZE_indelay,
	PLBPPCS1TATTRIBUTE  =>  PLBPPCS1TATTRIBUTE_indelay,
	PLBPPCS1TYPE  =>  PLBPPCS1TYPE_indelay,
	PLBPPCS1UABUS  =>  PLBPPCS1UABUS_indelay,
	PLBPPCS1WRBURST  =>  PLBPPCS1WRBURST_indelay,
	PLBPPCS1WRDBUS  =>  PLBPPCS1WRDBUS_indelay,
	PLBPPCS1WRPENDPRI  =>  PLBPPCS1WRPENDPRI_indelay,
	PLBPPCS1WRPENDREQ  =>  PLBPPCS1WRPENDREQ_indelay,
	PLBPPCS1WRPRIM  =>  PLBPPCS1WRPRIM_indelay,
	RSTC440RESETCHIP  =>  RSTC440RESETCHIP_indelay,
	RSTC440RESETCORE  =>  RSTC440RESETCORE_indelay,
	RSTC440RESETSYSTEM  =>  RSTC440RESETSYSTEM_indelay,
	TIEC440DCURDLDCACHEPLBPRIO  =>  TIEC440DCURDLDCACHEPLBPRIO_indelay,
	TIEC440DCURDNONCACHEPLBPRIO  =>  TIEC440DCURDNONCACHEPLBPRIO_indelay,
	TIEC440DCURDTOUCHPLBPRIO  =>  TIEC440DCURDTOUCHPLBPRIO_indelay,
	TIEC440DCURDURGENTPLBPRIO  =>  TIEC440DCURDURGENTPLBPRIO_indelay,
	TIEC440DCUWRFLUSHPLBPRIO  =>  TIEC440DCUWRFLUSHPLBPRIO_indelay,
	TIEC440DCUWRSTOREPLBPRIO  =>  TIEC440DCUWRSTOREPLBPRIO_indelay,
	TIEC440DCUWRURGENTPLBPRIO  =>  TIEC440DCUWRURGENTPLBPRIO_indelay,
	TIEC440ENDIANRESET  =>  TIEC440ENDIANRESET_indelay,
	TIEC440ERPNRESET  =>  TIEC440ERPNRESET_indelay,
	TIEC440ICURDFETCHPLBPRIO  =>  TIEC440ICURDFETCHPLBPRIO_indelay,
	TIEC440ICURDSPECPLBPRIO  =>  TIEC440ICURDSPECPLBPRIO_indelay,
	TIEC440ICURDTOUCHPLBPRIO  =>  TIEC440ICURDTOUCHPLBPRIO_indelay,
	TIEC440PIR  =>  TIEC440PIR_indelay,
	TIEC440PVR  =>  TIEC440PVR_indelay,
	TIEC440USERRESET  =>  TIEC440USERRESET_indelay,
	TIEDCRBASEADDR  =>  TIEDCRBASEADDR_indelay,
	TRCC440TRACEDISABLE  =>  TRCC440TRACEDISABLE_indelay,
	TRCC440TRIGGEREVENTIN  =>  TRCC440TRIGGEREVENTIN_indelay
	);

	INIPROC : process
	begin
       case PPCS0_WIDTH_128N64 is
           when FALSE   =>  PPCS0_WIDTH_128N64_BINARY <= '0';
           when TRUE    =>  PPCS0_WIDTH_128N64_BINARY <= '1';
           when others  =>  assert FALSE report "Error : PPCS0_WIDTH_128N64 is neither TRUE nor FALSE." severity error;
       end case;
       case PPCS1_WIDTH_128N64 is
           when FALSE   =>  PPCS1_WIDTH_128N64_BINARY <= '0';
           when TRUE    =>  PPCS1_WIDTH_128N64_BINARY <= '1';
           when others  =>  assert FALSE report "Error : PPCS1_WIDTH_128N64 is neither TRUE nor FALSE." severity error;
       end case;
       case PPCDM_ASYNCMODE is
           when FALSE   =>  PPCDM_ASYNCMODE_BINARY <= '0';
           when TRUE    =>  PPCDM_ASYNCMODE_BINARY <= '1';
           when others  =>  assert FALSE report "Error : PPCDM_ASYNCMODE is neither TRUE nor FALSE." severity error;
       end case;
       case PPCDS_ASYNCMODE is
           when FALSE   =>  PPCDS_ASYNCMODE_BINARY <= '0';
           when TRUE    =>  PPCDS_ASYNCMODE_BINARY <= '1';
           when others  =>  assert FALSE report "Error : PPCDS_ASYNCMODE is neither TRUE nor FALSE." severity error;
       end case;
       case DCR_AUTOLOCK_ENABLE is
           when FALSE   =>  DCR_AUTOLOCK_ENABLE_BINARY <= '0';
           when TRUE    =>  DCR_AUTOLOCK_ENABLE_BINARY <= '1';
           when others  =>  assert FALSE report "Error : DCR_AUTOLOCK_ENABLE is neither TRUE nor FALSE." severity error;
       end case;
       case CLOCK_DELAY is
           when FALSE   =>  CLOCK_DELAY_BINARY <= "10000";
           when TRUE    =>  CLOCK_DELAY_BINARY <= "00000";
           when others  =>  assert FALSE report "Error : CLOCK_DELAY is neither TRUE nor FALSE." severity error;
       end case;
	wait;
	end process INIPROC;

	TIMING : process



	variable  DMA0LLRSTENGINEACK_GlitchData : VitalGlitchDataType;
	variable  DMA0LLRXDSTRDYN_GlitchData : VitalGlitchDataType;
	variable  DMA0LLTXD0_GlitchData : VitalGlitchDataType;
	variable  DMA0LLTXD1_GlitchData : VitalGlitchDataType;
	variable  DMA0LLTXD2_GlitchData : VitalGlitchDataType;
	variable  DMA0LLTXD3_GlitchData : VitalGlitchDataType;
	variable  DMA0LLTXD4_GlitchData : VitalGlitchDataType;
	variable  DMA0LLTXD5_GlitchData : VitalGlitchDataType;
	variable  DMA0LLTXD6_GlitchData : VitalGlitchDataType;
	variable  DMA0LLTXD7_GlitchData : VitalGlitchDataType;
	variable  DMA0LLTXD8_GlitchData : VitalGlitchDataType;
	variable  DMA0LLTXD9_GlitchData : VitalGlitchDataType;
	variable  DMA0LLTXD10_GlitchData : VitalGlitchDataType;
	variable  DMA0LLTXD11_GlitchData : VitalGlitchDataType;
	variable  DMA0LLTXD12_GlitchData : VitalGlitchDataType;
	variable  DMA0LLTXD13_GlitchData : VitalGlitchDataType;
	variable  DMA0LLTXD14_GlitchData : VitalGlitchDataType;
	variable  DMA0LLTXD15_GlitchData : VitalGlitchDataType;
	variable  DMA0LLTXD16_GlitchData : VitalGlitchDataType;
	variable  DMA0LLTXD17_GlitchData : VitalGlitchDataType;
	variable  DMA0LLTXD18_GlitchData : VitalGlitchDataType;
	variable  DMA0LLTXD19_GlitchData : VitalGlitchDataType;
	variable  DMA0LLTXD20_GlitchData : VitalGlitchDataType;
	variable  DMA0LLTXD21_GlitchData : VitalGlitchDataType;
	variable  DMA0LLTXD22_GlitchData : VitalGlitchDataType;
	variable  DMA0LLTXD23_GlitchData : VitalGlitchDataType;
	variable  DMA0LLTXD24_GlitchData : VitalGlitchDataType;
	variable  DMA0LLTXD25_GlitchData : VitalGlitchDataType;
	variable  DMA0LLTXD26_GlitchData : VitalGlitchDataType;
	variable  DMA0LLTXD27_GlitchData : VitalGlitchDataType;
	variable  DMA0LLTXD28_GlitchData : VitalGlitchDataType;
	variable  DMA0LLTXD29_GlitchData : VitalGlitchDataType;
	variable  DMA0LLTXD30_GlitchData : VitalGlitchDataType;
	variable  DMA0LLTXD31_GlitchData : VitalGlitchDataType;
	variable  DMA0LLTXEOFN_GlitchData : VitalGlitchDataType;
	variable  DMA0LLTXEOPN_GlitchData : VitalGlitchDataType;
	variable  DMA0LLTXREM0_GlitchData : VitalGlitchDataType;
	variable  DMA0LLTXREM1_GlitchData : VitalGlitchDataType;
	variable  DMA0LLTXREM2_GlitchData : VitalGlitchDataType;
	variable  DMA0LLTXREM3_GlitchData : VitalGlitchDataType;
	variable  DMA0LLTXSOFN_GlitchData : VitalGlitchDataType;
	variable  DMA0LLTXSOPN_GlitchData : VitalGlitchDataType;
	variable  DMA0LLTXSRCRDYN_GlitchData : VitalGlitchDataType;
	variable  DMA0RXIRQ_GlitchData : VitalGlitchDataType;
	variable  DMA0TXIRQ_GlitchData : VitalGlitchDataType;
	variable  DMA1LLRSTENGINEACK_GlitchData : VitalGlitchDataType;
	variable  DMA1LLRXDSTRDYN_GlitchData : VitalGlitchDataType;
	variable  DMA1LLTXD0_GlitchData : VitalGlitchDataType;
	variable  DMA1LLTXD1_GlitchData : VitalGlitchDataType;
	variable  DMA1LLTXD2_GlitchData : VitalGlitchDataType;
	variable  DMA1LLTXD3_GlitchData : VitalGlitchDataType;
	variable  DMA1LLTXD4_GlitchData : VitalGlitchDataType;
	variable  DMA1LLTXD5_GlitchData : VitalGlitchDataType;
	variable  DMA1LLTXD6_GlitchData : VitalGlitchDataType;
	variable  DMA1LLTXD7_GlitchData : VitalGlitchDataType;
	variable  DMA1LLTXD8_GlitchData : VitalGlitchDataType;
	variable  DMA1LLTXD9_GlitchData : VitalGlitchDataType;
	variable  DMA1LLTXD10_GlitchData : VitalGlitchDataType;
	variable  DMA1LLTXD11_GlitchData : VitalGlitchDataType;
	variable  DMA1LLTXD12_GlitchData : VitalGlitchDataType;
	variable  DMA1LLTXD13_GlitchData : VitalGlitchDataType;
	variable  DMA1LLTXD14_GlitchData : VitalGlitchDataType;
	variable  DMA1LLTXD15_GlitchData : VitalGlitchDataType;
	variable  DMA1LLTXD16_GlitchData : VitalGlitchDataType;
	variable  DMA1LLTXD17_GlitchData : VitalGlitchDataType;
	variable  DMA1LLTXD18_GlitchData : VitalGlitchDataType;
	variable  DMA1LLTXD19_GlitchData : VitalGlitchDataType;
	variable  DMA1LLTXD20_GlitchData : VitalGlitchDataType;
	variable  DMA1LLTXD21_GlitchData : VitalGlitchDataType;
	variable  DMA1LLTXD22_GlitchData : VitalGlitchDataType;
	variable  DMA1LLTXD23_GlitchData : VitalGlitchDataType;
	variable  DMA1LLTXD24_GlitchData : VitalGlitchDataType;
	variable  DMA1LLTXD25_GlitchData : VitalGlitchDataType;
	variable  DMA1LLTXD26_GlitchData : VitalGlitchDataType;
	variable  DMA1LLTXD27_GlitchData : VitalGlitchDataType;
	variable  DMA1LLTXD28_GlitchData : VitalGlitchDataType;
	variable  DMA1LLTXD29_GlitchData : VitalGlitchDataType;
	variable  DMA1LLTXD30_GlitchData : VitalGlitchDataType;
	variable  DMA1LLTXD31_GlitchData : VitalGlitchDataType;
	variable  DMA1LLTXEOFN_GlitchData : VitalGlitchDataType;
	variable  DMA1LLTXEOPN_GlitchData : VitalGlitchDataType;
	variable  DMA1LLTXREM0_GlitchData : VitalGlitchDataType;
	variable  DMA1LLTXREM1_GlitchData : VitalGlitchDataType;
	variable  DMA1LLTXREM2_GlitchData : VitalGlitchDataType;
	variable  DMA1LLTXREM3_GlitchData : VitalGlitchDataType;
	variable  DMA1LLTXSOFN_GlitchData : VitalGlitchDataType;
	variable  DMA1LLTXSOPN_GlitchData : VitalGlitchDataType;
	variable  DMA1LLTXSRCRDYN_GlitchData : VitalGlitchDataType;
	variable  DMA1RXIRQ_GlitchData : VitalGlitchDataType;
	variable  DMA1TXIRQ_GlitchData : VitalGlitchDataType;
	variable  DMA2LLRSTENGINEACK_GlitchData : VitalGlitchDataType;
	variable  DMA2LLRXDSTRDYN_GlitchData : VitalGlitchDataType;
	variable  DMA2LLTXD0_GlitchData : VitalGlitchDataType;
	variable  DMA2LLTXD1_GlitchData : VitalGlitchDataType;
	variable  DMA2LLTXD2_GlitchData : VitalGlitchDataType;
	variable  DMA2LLTXD3_GlitchData : VitalGlitchDataType;
	variable  DMA2LLTXD4_GlitchData : VitalGlitchDataType;
	variable  DMA2LLTXD5_GlitchData : VitalGlitchDataType;
	variable  DMA2LLTXD6_GlitchData : VitalGlitchDataType;
	variable  DMA2LLTXD7_GlitchData : VitalGlitchDataType;
	variable  DMA2LLTXD8_GlitchData : VitalGlitchDataType;
	variable  DMA2LLTXD9_GlitchData : VitalGlitchDataType;
	variable  DMA2LLTXD10_GlitchData : VitalGlitchDataType;
	variable  DMA2LLTXD11_GlitchData : VitalGlitchDataType;
	variable  DMA2LLTXD12_GlitchData : VitalGlitchDataType;
	variable  DMA2LLTXD13_GlitchData : VitalGlitchDataType;
	variable  DMA2LLTXD14_GlitchData : VitalGlitchDataType;
	variable  DMA2LLTXD15_GlitchData : VitalGlitchDataType;
	variable  DMA2LLTXD16_GlitchData : VitalGlitchDataType;
	variable  DMA2LLTXD17_GlitchData : VitalGlitchDataType;
	variable  DMA2LLTXD18_GlitchData : VitalGlitchDataType;
	variable  DMA2LLTXD19_GlitchData : VitalGlitchDataType;
	variable  DMA2LLTXD20_GlitchData : VitalGlitchDataType;
	variable  DMA2LLTXD21_GlitchData : VitalGlitchDataType;
	variable  DMA2LLTXD22_GlitchData : VitalGlitchDataType;
	variable  DMA2LLTXD23_GlitchData : VitalGlitchDataType;
	variable  DMA2LLTXD24_GlitchData : VitalGlitchDataType;
	variable  DMA2LLTXD25_GlitchData : VitalGlitchDataType;
	variable  DMA2LLTXD26_GlitchData : VitalGlitchDataType;
	variable  DMA2LLTXD27_GlitchData : VitalGlitchDataType;
	variable  DMA2LLTXD28_GlitchData : VitalGlitchDataType;
	variable  DMA2LLTXD29_GlitchData : VitalGlitchDataType;
	variable  DMA2LLTXD30_GlitchData : VitalGlitchDataType;
	variable  DMA2LLTXD31_GlitchData : VitalGlitchDataType;
	variable  DMA2LLTXEOFN_GlitchData : VitalGlitchDataType;
	variable  DMA2LLTXEOPN_GlitchData : VitalGlitchDataType;
	variable  DMA2LLTXREM0_GlitchData : VitalGlitchDataType;
	variable  DMA2LLTXREM1_GlitchData : VitalGlitchDataType;
	variable  DMA2LLTXREM2_GlitchData : VitalGlitchDataType;
	variable  DMA2LLTXREM3_GlitchData : VitalGlitchDataType;
	variable  DMA2LLTXSOFN_GlitchData : VitalGlitchDataType;
	variable  DMA2LLTXSOPN_GlitchData : VitalGlitchDataType;
	variable  DMA2LLTXSRCRDYN_GlitchData : VitalGlitchDataType;
	variable  DMA2RXIRQ_GlitchData : VitalGlitchDataType;
	variable  DMA2TXIRQ_GlitchData : VitalGlitchDataType;
	variable  DMA3LLRSTENGINEACK_GlitchData : VitalGlitchDataType;
	variable  DMA3LLRXDSTRDYN_GlitchData : VitalGlitchDataType;
	variable  DMA3LLTXD0_GlitchData : VitalGlitchDataType;
	variable  DMA3LLTXD1_GlitchData : VitalGlitchDataType;
	variable  DMA3LLTXD2_GlitchData : VitalGlitchDataType;
	variable  DMA3LLTXD3_GlitchData : VitalGlitchDataType;
	variable  DMA3LLTXD4_GlitchData : VitalGlitchDataType;
	variable  DMA3LLTXD5_GlitchData : VitalGlitchDataType;
	variable  DMA3LLTXD6_GlitchData : VitalGlitchDataType;
	variable  DMA3LLTXD7_GlitchData : VitalGlitchDataType;
	variable  DMA3LLTXD8_GlitchData : VitalGlitchDataType;
	variable  DMA3LLTXD9_GlitchData : VitalGlitchDataType;
	variable  DMA3LLTXD10_GlitchData : VitalGlitchDataType;
	variable  DMA3LLTXD11_GlitchData : VitalGlitchDataType;
	variable  DMA3LLTXD12_GlitchData : VitalGlitchDataType;
	variable  DMA3LLTXD13_GlitchData : VitalGlitchDataType;
	variable  DMA3LLTXD14_GlitchData : VitalGlitchDataType;
	variable  DMA3LLTXD15_GlitchData : VitalGlitchDataType;
	variable  DMA3LLTXD16_GlitchData : VitalGlitchDataType;
	variable  DMA3LLTXD17_GlitchData : VitalGlitchDataType;
	variable  DMA3LLTXD18_GlitchData : VitalGlitchDataType;
	variable  DMA3LLTXD19_GlitchData : VitalGlitchDataType;
	variable  DMA3LLTXD20_GlitchData : VitalGlitchDataType;
	variable  DMA3LLTXD21_GlitchData : VitalGlitchDataType;
	variable  DMA3LLTXD22_GlitchData : VitalGlitchDataType;
	variable  DMA3LLTXD23_GlitchData : VitalGlitchDataType;
	variable  DMA3LLTXD24_GlitchData : VitalGlitchDataType;
	variable  DMA3LLTXD25_GlitchData : VitalGlitchDataType;
	variable  DMA3LLTXD26_GlitchData : VitalGlitchDataType;
	variable  DMA3LLTXD27_GlitchData : VitalGlitchDataType;
	variable  DMA3LLTXD28_GlitchData : VitalGlitchDataType;
	variable  DMA3LLTXD29_GlitchData : VitalGlitchDataType;
	variable  DMA3LLTXD30_GlitchData : VitalGlitchDataType;
	variable  DMA3LLTXD31_GlitchData : VitalGlitchDataType;
	variable  DMA3LLTXEOFN_GlitchData : VitalGlitchDataType;
	variable  DMA3LLTXEOPN_GlitchData : VitalGlitchDataType;
	variable  DMA3LLTXREM0_GlitchData : VitalGlitchDataType;
	variable  DMA3LLTXREM1_GlitchData : VitalGlitchDataType;
	variable  DMA3LLTXREM2_GlitchData : VitalGlitchDataType;
	variable  DMA3LLTXREM3_GlitchData : VitalGlitchDataType;
	variable  DMA3LLTXSOFN_GlitchData : VitalGlitchDataType;
	variable  DMA3LLTXSOPN_GlitchData : VitalGlitchDataType;
	variable  DMA3LLTXSRCRDYN_GlitchData : VitalGlitchDataType;
	variable  DMA3RXIRQ_GlitchData : VitalGlitchDataType;
	variable  DMA3TXIRQ_GlitchData : VitalGlitchDataType;
	variable  PPCDMDCRABUS0_GlitchData : VitalGlitchDataType;
	variable  PPCDMDCRABUS1_GlitchData : VitalGlitchDataType;
	variable  PPCDMDCRABUS2_GlitchData : VitalGlitchDataType;
	variable  PPCDMDCRABUS3_GlitchData : VitalGlitchDataType;
	variable  PPCDMDCRABUS4_GlitchData : VitalGlitchDataType;
	variable  PPCDMDCRABUS5_GlitchData : VitalGlitchDataType;
	variable  PPCDMDCRABUS6_GlitchData : VitalGlitchDataType;
	variable  PPCDMDCRABUS7_GlitchData : VitalGlitchDataType;
	variable  PPCDMDCRABUS8_GlitchData : VitalGlitchDataType;
	variable  PPCDMDCRABUS9_GlitchData : VitalGlitchDataType;
	variable  PPCDMDCRDBUSOUT0_GlitchData : VitalGlitchDataType;
	variable  PPCDMDCRDBUSOUT1_GlitchData : VitalGlitchDataType;
	variable  PPCDMDCRDBUSOUT2_GlitchData : VitalGlitchDataType;
	variable  PPCDMDCRDBUSOUT3_GlitchData : VitalGlitchDataType;
	variable  PPCDMDCRDBUSOUT4_GlitchData : VitalGlitchDataType;
	variable  PPCDMDCRDBUSOUT5_GlitchData : VitalGlitchDataType;
	variable  PPCDMDCRDBUSOUT6_GlitchData : VitalGlitchDataType;
	variable  PPCDMDCRDBUSOUT7_GlitchData : VitalGlitchDataType;
	variable  PPCDMDCRDBUSOUT8_GlitchData : VitalGlitchDataType;
	variable  PPCDMDCRDBUSOUT9_GlitchData : VitalGlitchDataType;
	variable  PPCDMDCRDBUSOUT10_GlitchData : VitalGlitchDataType;
	variable  PPCDMDCRDBUSOUT11_GlitchData : VitalGlitchDataType;
	variable  PPCDMDCRDBUSOUT12_GlitchData : VitalGlitchDataType;
	variable  PPCDMDCRDBUSOUT13_GlitchData : VitalGlitchDataType;
	variable  PPCDMDCRDBUSOUT14_GlitchData : VitalGlitchDataType;
	variable  PPCDMDCRDBUSOUT15_GlitchData : VitalGlitchDataType;
	variable  PPCDMDCRDBUSOUT16_GlitchData : VitalGlitchDataType;
	variable  PPCDMDCRDBUSOUT17_GlitchData : VitalGlitchDataType;
	variable  PPCDMDCRDBUSOUT18_GlitchData : VitalGlitchDataType;
	variable  PPCDMDCRDBUSOUT19_GlitchData : VitalGlitchDataType;
	variable  PPCDMDCRDBUSOUT20_GlitchData : VitalGlitchDataType;
	variable  PPCDMDCRDBUSOUT21_GlitchData : VitalGlitchDataType;
	variable  PPCDMDCRDBUSOUT22_GlitchData : VitalGlitchDataType;
	variable  PPCDMDCRDBUSOUT23_GlitchData : VitalGlitchDataType;
	variable  PPCDMDCRDBUSOUT24_GlitchData : VitalGlitchDataType;
	variable  PPCDMDCRDBUSOUT25_GlitchData : VitalGlitchDataType;
	variable  PPCDMDCRDBUSOUT26_GlitchData : VitalGlitchDataType;
	variable  PPCDMDCRDBUSOUT27_GlitchData : VitalGlitchDataType;
	variable  PPCDMDCRDBUSOUT28_GlitchData : VitalGlitchDataType;
	variable  PPCDMDCRDBUSOUT29_GlitchData : VitalGlitchDataType;
	variable  PPCDMDCRDBUSOUT30_GlitchData : VitalGlitchDataType;
	variable  PPCDMDCRDBUSOUT31_GlitchData : VitalGlitchDataType;
	variable  PPCDMDCRREAD_GlitchData : VitalGlitchDataType;
	variable  PPCDMDCRUABUS20_GlitchData : VitalGlitchDataType;
	variable  PPCDMDCRUABUS21_GlitchData : VitalGlitchDataType;
	variable  PPCDMDCRWRITE_GlitchData : VitalGlitchDataType;
	variable  PPCMPLBABORT_GlitchData : VitalGlitchDataType;
	variable  PPCMPLBABUS0_GlitchData : VitalGlitchDataType;
	variable  PPCMPLBABUS1_GlitchData : VitalGlitchDataType;
	variable  PPCMPLBABUS2_GlitchData : VitalGlitchDataType;
	variable  PPCMPLBABUS3_GlitchData : VitalGlitchDataType;
	variable  PPCMPLBABUS4_GlitchData : VitalGlitchDataType;
	variable  PPCMPLBABUS5_GlitchData : VitalGlitchDataType;
	variable  PPCMPLBABUS6_GlitchData : VitalGlitchDataType;
	variable  PPCMPLBABUS7_GlitchData : VitalGlitchDataType;
	variable  PPCMPLBABUS8_GlitchData : VitalGlitchDataType;
	variable  PPCMPLBABUS9_GlitchData : VitalGlitchDataType;
	variable  PPCMPLBABUS10_GlitchData : VitalGlitchDataType;
	variable  PPCMPLBABUS11_GlitchData : VitalGlitchDataType;
	variable  PPCMPLBABUS12_GlitchData : VitalGlitchDataType;
	variable  PPCMPLBABUS13_GlitchData : VitalGlitchDataType;
	variable  PPCMPLBABUS14_GlitchData : VitalGlitchDataType;
	variable  PPCMPLBABUS15_GlitchData : VitalGlitchDataType;
	variable  PPCMPLBABUS16_GlitchData : VitalGlitchDataType;
	variable  PPCMPLBABUS17_GlitchData : VitalGlitchDataType;
	variable  PPCMPLBABUS18_GlitchData : VitalGlitchDataType;
	variable  PPCMPLBABUS19_GlitchData : VitalGlitchDataType;
	variable  PPCMPLBABUS20_GlitchData : VitalGlitchDataType;
	variable  PPCMPLBABUS21_GlitchData : VitalGlitchDataType;
	variable  PPCMPLBABUS22_GlitchData : VitalGlitchDataType;
	variable  PPCMPLBABUS23_GlitchData : VitalGlitchDataType;
	variable  PPCMPLBABUS24_GlitchData : VitalGlitchDataType;
	variable  PPCMPLBABUS25_GlitchData : VitalGlitchDataType;
	variable  PPCMPLBABUS26_GlitchData : VitalGlitchDataType;
	variable  PPCMPLBABUS27_GlitchData : VitalGlitchDataType;
	variable  PPCMPLBABUS28_GlitchData : VitalGlitchDataType;
	variable  PPCMPLBABUS29_GlitchData : VitalGlitchDataType;
	variable  PPCMPLBABUS30_GlitchData : VitalGlitchDataType;
	variable  PPCMPLBABUS31_GlitchData : VitalGlitchDataType;
	variable  PPCMPLBBE0_GlitchData : VitalGlitchDataType;
	variable  PPCMPLBBE1_GlitchData : VitalGlitchDataType;
	variable  PPCMPLBBE2_GlitchData : VitalGlitchDataType;
	variable  PPCMPLBBE3_GlitchData : VitalGlitchDataType;
	variable  PPCMPLBBE4_GlitchData : VitalGlitchDataType;
	variable  PPCMPLBBE5_GlitchData : VitalGlitchDataType;
	variable  PPCMPLBBE6_GlitchData : VitalGlitchDataType;
	variable  PPCMPLBBE7_GlitchData : VitalGlitchDataType;
	variable  PPCMPLBBE8_GlitchData : VitalGlitchDataType;
	variable  PPCMPLBBE9_GlitchData : VitalGlitchDataType;
	variable  PPCMPLBBE10_GlitchData : VitalGlitchDataType;
	variable  PPCMPLBBE11_GlitchData : VitalGlitchDataType;
	variable  PPCMPLBBE12_GlitchData : VitalGlitchDataType;
	variable  PPCMPLBBE13_GlitchData : VitalGlitchDataType;
	variable  PPCMPLBBE14_GlitchData : VitalGlitchDataType;
	variable  PPCMPLBBE15_GlitchData : VitalGlitchDataType;
	variable  PPCMPLBBUSLOCK_GlitchData : VitalGlitchDataType;
	variable  PPCMPLBLOCKERR_GlitchData : VitalGlitchDataType;
	variable  PPCMPLBPRIORITY0_GlitchData : VitalGlitchDataType;
	variable  PPCMPLBPRIORITY1_GlitchData : VitalGlitchDataType;
	variable  PPCMPLBRDBURST_GlitchData : VitalGlitchDataType;
	variable  PPCMPLBREQUEST_GlitchData : VitalGlitchDataType;
	variable  PPCMPLBRNW_GlitchData : VitalGlitchDataType;
	variable  PPCMPLBSIZE0_GlitchData : VitalGlitchDataType;
	variable  PPCMPLBSIZE1_GlitchData : VitalGlitchDataType;
	variable  PPCMPLBSIZE2_GlitchData : VitalGlitchDataType;
	variable  PPCMPLBSIZE3_GlitchData : VitalGlitchDataType;
	variable  PPCMPLBTATTRIBUTE0_GlitchData : VitalGlitchDataType;
	variable  PPCMPLBTATTRIBUTE1_GlitchData : VitalGlitchDataType;
	variable  PPCMPLBTATTRIBUTE2_GlitchData : VitalGlitchDataType;
	variable  PPCMPLBTATTRIBUTE3_GlitchData : VitalGlitchDataType;
	variable  PPCMPLBTATTRIBUTE4_GlitchData : VitalGlitchDataType;
	variable  PPCMPLBTATTRIBUTE5_GlitchData : VitalGlitchDataType;
	variable  PPCMPLBTATTRIBUTE6_GlitchData : VitalGlitchDataType;
	variable  PPCMPLBTATTRIBUTE7_GlitchData : VitalGlitchDataType;
	variable  PPCMPLBTATTRIBUTE8_GlitchData : VitalGlitchDataType;
	variable  PPCMPLBTATTRIBUTE9_GlitchData : VitalGlitchDataType;
	variable  PPCMPLBTATTRIBUTE10_GlitchData : VitalGlitchDataType;
	variable  PPCMPLBTATTRIBUTE11_GlitchData : VitalGlitchDataType;
	variable  PPCMPLBTATTRIBUTE12_GlitchData : VitalGlitchDataType;
	variable  PPCMPLBTATTRIBUTE13_GlitchData : VitalGlitchDataType;
	variable  PPCMPLBTATTRIBUTE14_GlitchData : VitalGlitchDataType;
	variable  PPCMPLBTATTRIBUTE15_GlitchData : VitalGlitchDataType;
	variable  PPCMPLBTYPE0_GlitchData : VitalGlitchDataType;
	variable  PPCMPLBTYPE1_GlitchData : VitalGlitchDataType;
	variable  PPCMPLBTYPE2_GlitchData : VitalGlitchDataType;
	variable  PPCMPLBUABUS28_GlitchData : VitalGlitchDataType;
	variable  PPCMPLBUABUS29_GlitchData : VitalGlitchDataType;
	variable  PPCMPLBUABUS30_GlitchData : VitalGlitchDataType;
	variable  PPCMPLBUABUS31_GlitchData : VitalGlitchDataType;
	variable  PPCMPLBWRBURST_GlitchData : VitalGlitchDataType;
	variable  PPCMPLBWRDBUS0_GlitchData : VitalGlitchDataType;
	variable  PPCMPLBWRDBUS1_GlitchData : VitalGlitchDataType;
	variable  PPCMPLBWRDBUS2_GlitchData : VitalGlitchDataType;
	variable  PPCMPLBWRDBUS3_GlitchData : VitalGlitchDataType;
	variable  PPCMPLBWRDBUS4_GlitchData : VitalGlitchDataType;
	variable  PPCMPLBWRDBUS5_GlitchData : VitalGlitchDataType;
	variable  PPCMPLBWRDBUS6_GlitchData : VitalGlitchDataType;
	variable  PPCMPLBWRDBUS7_GlitchData : VitalGlitchDataType;
	variable  PPCMPLBWRDBUS8_GlitchData : VitalGlitchDataType;
	variable  PPCMPLBWRDBUS9_GlitchData : VitalGlitchDataType;
	variable  PPCMPLBWRDBUS10_GlitchData : VitalGlitchDataType;
	variable  PPCMPLBWRDBUS11_GlitchData : VitalGlitchDataType;
	variable  PPCMPLBWRDBUS12_GlitchData : VitalGlitchDataType;
	variable  PPCMPLBWRDBUS13_GlitchData : VitalGlitchDataType;
	variable  PPCMPLBWRDBUS14_GlitchData : VitalGlitchDataType;
	variable  PPCMPLBWRDBUS15_GlitchData : VitalGlitchDataType;
	variable  PPCMPLBWRDBUS16_GlitchData : VitalGlitchDataType;
	variable  PPCMPLBWRDBUS17_GlitchData : VitalGlitchDataType;
	variable  PPCMPLBWRDBUS18_GlitchData : VitalGlitchDataType;
	variable  PPCMPLBWRDBUS19_GlitchData : VitalGlitchDataType;
	variable  PPCMPLBWRDBUS20_GlitchData : VitalGlitchDataType;
	variable  PPCMPLBWRDBUS21_GlitchData : VitalGlitchDataType;
	variable  PPCMPLBWRDBUS22_GlitchData : VitalGlitchDataType;
	variable  PPCMPLBWRDBUS23_GlitchData : VitalGlitchDataType;
	variable  PPCMPLBWRDBUS24_GlitchData : VitalGlitchDataType;
	variable  PPCMPLBWRDBUS25_GlitchData : VitalGlitchDataType;
	variable  PPCMPLBWRDBUS26_GlitchData : VitalGlitchDataType;
	variable  PPCMPLBWRDBUS27_GlitchData : VitalGlitchDataType;
	variable  PPCMPLBWRDBUS28_GlitchData : VitalGlitchDataType;
	variable  PPCMPLBWRDBUS29_GlitchData : VitalGlitchDataType;
	variable  PPCMPLBWRDBUS30_GlitchData : VitalGlitchDataType;
	variable  PPCMPLBWRDBUS31_GlitchData : VitalGlitchDataType;
	variable  PPCMPLBWRDBUS32_GlitchData : VitalGlitchDataType;
	variable  PPCMPLBWRDBUS33_GlitchData : VitalGlitchDataType;
	variable  PPCMPLBWRDBUS34_GlitchData : VitalGlitchDataType;
	variable  PPCMPLBWRDBUS35_GlitchData : VitalGlitchDataType;
	variable  PPCMPLBWRDBUS36_GlitchData : VitalGlitchDataType;
	variable  PPCMPLBWRDBUS37_GlitchData : VitalGlitchDataType;
	variable  PPCMPLBWRDBUS38_GlitchData : VitalGlitchDataType;
	variable  PPCMPLBWRDBUS39_GlitchData : VitalGlitchDataType;
	variable  PPCMPLBWRDBUS40_GlitchData : VitalGlitchDataType;
	variable  PPCMPLBWRDBUS41_GlitchData : VitalGlitchDataType;
	variable  PPCMPLBWRDBUS42_GlitchData : VitalGlitchDataType;
	variable  PPCMPLBWRDBUS43_GlitchData : VitalGlitchDataType;
	variable  PPCMPLBWRDBUS44_GlitchData : VitalGlitchDataType;
	variable  PPCMPLBWRDBUS45_GlitchData : VitalGlitchDataType;
	variable  PPCMPLBWRDBUS46_GlitchData : VitalGlitchDataType;
	variable  PPCMPLBWRDBUS47_GlitchData : VitalGlitchDataType;
	variable  PPCMPLBWRDBUS48_GlitchData : VitalGlitchDataType;
	variable  PPCMPLBWRDBUS49_GlitchData : VitalGlitchDataType;
	variable  PPCMPLBWRDBUS50_GlitchData : VitalGlitchDataType;
	variable  PPCMPLBWRDBUS51_GlitchData : VitalGlitchDataType;
	variable  PPCMPLBWRDBUS52_GlitchData : VitalGlitchDataType;
	variable  PPCMPLBWRDBUS53_GlitchData : VitalGlitchDataType;
	variable  PPCMPLBWRDBUS54_GlitchData : VitalGlitchDataType;
	variable  PPCMPLBWRDBUS55_GlitchData : VitalGlitchDataType;
	variable  PPCMPLBWRDBUS56_GlitchData : VitalGlitchDataType;
	variable  PPCMPLBWRDBUS57_GlitchData : VitalGlitchDataType;
	variable  PPCMPLBWRDBUS58_GlitchData : VitalGlitchDataType;
	variable  PPCMPLBWRDBUS59_GlitchData : VitalGlitchDataType;
	variable  PPCMPLBWRDBUS60_GlitchData : VitalGlitchDataType;
	variable  PPCMPLBWRDBUS61_GlitchData : VitalGlitchDataType;
	variable  PPCMPLBWRDBUS62_GlitchData : VitalGlitchDataType;
	variable  PPCMPLBWRDBUS63_GlitchData : VitalGlitchDataType;
	variable  PPCMPLBWRDBUS64_GlitchData : VitalGlitchDataType;
	variable  PPCMPLBWRDBUS65_GlitchData : VitalGlitchDataType;
	variable  PPCMPLBWRDBUS66_GlitchData : VitalGlitchDataType;
	variable  PPCMPLBWRDBUS67_GlitchData : VitalGlitchDataType;
	variable  PPCMPLBWRDBUS68_GlitchData : VitalGlitchDataType;
	variable  PPCMPLBWRDBUS69_GlitchData : VitalGlitchDataType;
	variable  PPCMPLBWRDBUS70_GlitchData : VitalGlitchDataType;
	variable  PPCMPLBWRDBUS71_GlitchData : VitalGlitchDataType;
	variable  PPCMPLBWRDBUS72_GlitchData : VitalGlitchDataType;
	variable  PPCMPLBWRDBUS73_GlitchData : VitalGlitchDataType;
	variable  PPCMPLBWRDBUS74_GlitchData : VitalGlitchDataType;
	variable  PPCMPLBWRDBUS75_GlitchData : VitalGlitchDataType;
	variable  PPCMPLBWRDBUS76_GlitchData : VitalGlitchDataType;
	variable  PPCMPLBWRDBUS77_GlitchData : VitalGlitchDataType;
	variable  PPCMPLBWRDBUS78_GlitchData : VitalGlitchDataType;
	variable  PPCMPLBWRDBUS79_GlitchData : VitalGlitchDataType;
	variable  PPCMPLBWRDBUS80_GlitchData : VitalGlitchDataType;
	variable  PPCMPLBWRDBUS81_GlitchData : VitalGlitchDataType;
	variable  PPCMPLBWRDBUS82_GlitchData : VitalGlitchDataType;
	variable  PPCMPLBWRDBUS83_GlitchData : VitalGlitchDataType;
	variable  PPCMPLBWRDBUS84_GlitchData : VitalGlitchDataType;
	variable  PPCMPLBWRDBUS85_GlitchData : VitalGlitchDataType;
	variable  PPCMPLBWRDBUS86_GlitchData : VitalGlitchDataType;
	variable  PPCMPLBWRDBUS87_GlitchData : VitalGlitchDataType;
	variable  PPCMPLBWRDBUS88_GlitchData : VitalGlitchDataType;
	variable  PPCMPLBWRDBUS89_GlitchData : VitalGlitchDataType;
	variable  PPCMPLBWRDBUS90_GlitchData : VitalGlitchDataType;
	variable  PPCMPLBWRDBUS91_GlitchData : VitalGlitchDataType;
	variable  PPCMPLBWRDBUS92_GlitchData : VitalGlitchDataType;
	variable  PPCMPLBWRDBUS93_GlitchData : VitalGlitchDataType;
	variable  PPCMPLBWRDBUS94_GlitchData : VitalGlitchDataType;
	variable  PPCMPLBWRDBUS95_GlitchData : VitalGlitchDataType;
	variable  PPCMPLBWRDBUS96_GlitchData : VitalGlitchDataType;
	variable  PPCMPLBWRDBUS97_GlitchData : VitalGlitchDataType;
	variable  PPCMPLBWRDBUS98_GlitchData : VitalGlitchDataType;
	variable  PPCMPLBWRDBUS99_GlitchData : VitalGlitchDataType;
	variable  PPCMPLBWRDBUS100_GlitchData : VitalGlitchDataType;
	variable  PPCMPLBWRDBUS101_GlitchData : VitalGlitchDataType;
	variable  PPCMPLBWRDBUS102_GlitchData : VitalGlitchDataType;
	variable  PPCMPLBWRDBUS103_GlitchData : VitalGlitchDataType;
	variable  PPCMPLBWRDBUS104_GlitchData : VitalGlitchDataType;
	variable  PPCMPLBWRDBUS105_GlitchData : VitalGlitchDataType;
	variable  PPCMPLBWRDBUS106_GlitchData : VitalGlitchDataType;
	variable  PPCMPLBWRDBUS107_GlitchData : VitalGlitchDataType;
	variable  PPCMPLBWRDBUS108_GlitchData : VitalGlitchDataType;
	variable  PPCMPLBWRDBUS109_GlitchData : VitalGlitchDataType;
	variable  PPCMPLBWRDBUS110_GlitchData : VitalGlitchDataType;
	variable  PPCMPLBWRDBUS111_GlitchData : VitalGlitchDataType;
	variable  PPCMPLBWRDBUS112_GlitchData : VitalGlitchDataType;
	variable  PPCMPLBWRDBUS113_GlitchData : VitalGlitchDataType;
	variable  PPCMPLBWRDBUS114_GlitchData : VitalGlitchDataType;
	variable  PPCMPLBWRDBUS115_GlitchData : VitalGlitchDataType;
	variable  PPCMPLBWRDBUS116_GlitchData : VitalGlitchDataType;
	variable  PPCMPLBWRDBUS117_GlitchData : VitalGlitchDataType;
	variable  PPCMPLBWRDBUS118_GlitchData : VitalGlitchDataType;
	variable  PPCMPLBWRDBUS119_GlitchData : VitalGlitchDataType;
	variable  PPCMPLBWRDBUS120_GlitchData : VitalGlitchDataType;
	variable  PPCMPLBWRDBUS121_GlitchData : VitalGlitchDataType;
	variable  PPCMPLBWRDBUS122_GlitchData : VitalGlitchDataType;
	variable  PPCMPLBWRDBUS123_GlitchData : VitalGlitchDataType;
	variable  PPCMPLBWRDBUS124_GlitchData : VitalGlitchDataType;
	variable  PPCMPLBWRDBUS125_GlitchData : VitalGlitchDataType;
	variable  PPCMPLBWRDBUS126_GlitchData : VitalGlitchDataType;
	variable  PPCMPLBWRDBUS127_GlitchData : VitalGlitchDataType;
	variable  PPCS0PLBADDRACK_GlitchData : VitalGlitchDataType;
	variable  PPCS0PLBMBUSY0_GlitchData : VitalGlitchDataType;
	variable  PPCS0PLBMBUSY1_GlitchData : VitalGlitchDataType;
	variable  PPCS0PLBMBUSY2_GlitchData : VitalGlitchDataType;
	variable  PPCS0PLBMBUSY3_GlitchData : VitalGlitchDataType;
	variable  PPCS0PLBMIRQ0_GlitchData : VitalGlitchDataType;
	variable  PPCS0PLBMIRQ1_GlitchData : VitalGlitchDataType;
	variable  PPCS0PLBMIRQ2_GlitchData : VitalGlitchDataType;
	variable  PPCS0PLBMIRQ3_GlitchData : VitalGlitchDataType;
	variable  PPCS0PLBMRDERR0_GlitchData : VitalGlitchDataType;
	variable  PPCS0PLBMRDERR1_GlitchData : VitalGlitchDataType;
	variable  PPCS0PLBMRDERR2_GlitchData : VitalGlitchDataType;
	variable  PPCS0PLBMRDERR3_GlitchData : VitalGlitchDataType;
	variable  PPCS0PLBMWRERR0_GlitchData : VitalGlitchDataType;
	variable  PPCS0PLBMWRERR1_GlitchData : VitalGlitchDataType;
	variable  PPCS0PLBMWRERR2_GlitchData : VitalGlitchDataType;
	variable  PPCS0PLBMWRERR3_GlitchData : VitalGlitchDataType;
	variable  PPCS0PLBRDBTERM_GlitchData : VitalGlitchDataType;
	variable  PPCS0PLBRDCOMP_GlitchData : VitalGlitchDataType;
	variable  PPCS0PLBRDDACK_GlitchData : VitalGlitchDataType;
	variable  PPCS0PLBRDDBUS0_GlitchData : VitalGlitchDataType;
	variable  PPCS0PLBRDDBUS1_GlitchData : VitalGlitchDataType;
	variable  PPCS0PLBRDDBUS2_GlitchData : VitalGlitchDataType;
	variable  PPCS0PLBRDDBUS3_GlitchData : VitalGlitchDataType;
	variable  PPCS0PLBRDDBUS4_GlitchData : VitalGlitchDataType;
	variable  PPCS0PLBRDDBUS5_GlitchData : VitalGlitchDataType;
	variable  PPCS0PLBRDDBUS6_GlitchData : VitalGlitchDataType;
	variable  PPCS0PLBRDDBUS7_GlitchData : VitalGlitchDataType;
	variable  PPCS0PLBRDDBUS8_GlitchData : VitalGlitchDataType;
	variable  PPCS0PLBRDDBUS9_GlitchData : VitalGlitchDataType;
	variable  PPCS0PLBRDDBUS10_GlitchData : VitalGlitchDataType;
	variable  PPCS0PLBRDDBUS11_GlitchData : VitalGlitchDataType;
	variable  PPCS0PLBRDDBUS12_GlitchData : VitalGlitchDataType;
	variable  PPCS0PLBRDDBUS13_GlitchData : VitalGlitchDataType;
	variable  PPCS0PLBRDDBUS14_GlitchData : VitalGlitchDataType;
	variable  PPCS0PLBRDDBUS15_GlitchData : VitalGlitchDataType;
	variable  PPCS0PLBRDDBUS16_GlitchData : VitalGlitchDataType;
	variable  PPCS0PLBRDDBUS17_GlitchData : VitalGlitchDataType;
	variable  PPCS0PLBRDDBUS18_GlitchData : VitalGlitchDataType;
	variable  PPCS0PLBRDDBUS19_GlitchData : VitalGlitchDataType;
	variable  PPCS0PLBRDDBUS20_GlitchData : VitalGlitchDataType;
	variable  PPCS0PLBRDDBUS21_GlitchData : VitalGlitchDataType;
	variable  PPCS0PLBRDDBUS22_GlitchData : VitalGlitchDataType;
	variable  PPCS0PLBRDDBUS23_GlitchData : VitalGlitchDataType;
	variable  PPCS0PLBRDDBUS24_GlitchData : VitalGlitchDataType;
	variable  PPCS0PLBRDDBUS25_GlitchData : VitalGlitchDataType;
	variable  PPCS0PLBRDDBUS26_GlitchData : VitalGlitchDataType;
	variable  PPCS0PLBRDDBUS27_GlitchData : VitalGlitchDataType;
	variable  PPCS0PLBRDDBUS28_GlitchData : VitalGlitchDataType;
	variable  PPCS0PLBRDDBUS29_GlitchData : VitalGlitchDataType;
	variable  PPCS0PLBRDDBUS30_GlitchData : VitalGlitchDataType;
	variable  PPCS0PLBRDDBUS31_GlitchData : VitalGlitchDataType;
	variable  PPCS0PLBRDDBUS32_GlitchData : VitalGlitchDataType;
	variable  PPCS0PLBRDDBUS33_GlitchData : VitalGlitchDataType;
	variable  PPCS0PLBRDDBUS34_GlitchData : VitalGlitchDataType;
	variable  PPCS0PLBRDDBUS35_GlitchData : VitalGlitchDataType;
	variable  PPCS0PLBRDDBUS36_GlitchData : VitalGlitchDataType;
	variable  PPCS0PLBRDDBUS37_GlitchData : VitalGlitchDataType;
	variable  PPCS0PLBRDDBUS38_GlitchData : VitalGlitchDataType;
	variable  PPCS0PLBRDDBUS39_GlitchData : VitalGlitchDataType;
	variable  PPCS0PLBRDDBUS40_GlitchData : VitalGlitchDataType;
	variable  PPCS0PLBRDDBUS41_GlitchData : VitalGlitchDataType;
	variable  PPCS0PLBRDDBUS42_GlitchData : VitalGlitchDataType;
	variable  PPCS0PLBRDDBUS43_GlitchData : VitalGlitchDataType;
	variable  PPCS0PLBRDDBUS44_GlitchData : VitalGlitchDataType;
	variable  PPCS0PLBRDDBUS45_GlitchData : VitalGlitchDataType;
	variable  PPCS0PLBRDDBUS46_GlitchData : VitalGlitchDataType;
	variable  PPCS0PLBRDDBUS47_GlitchData : VitalGlitchDataType;
	variable  PPCS0PLBRDDBUS48_GlitchData : VitalGlitchDataType;
	variable  PPCS0PLBRDDBUS49_GlitchData : VitalGlitchDataType;
	variable  PPCS0PLBRDDBUS50_GlitchData : VitalGlitchDataType;
	variable  PPCS0PLBRDDBUS51_GlitchData : VitalGlitchDataType;
	variable  PPCS0PLBRDDBUS52_GlitchData : VitalGlitchDataType;
	variable  PPCS0PLBRDDBUS53_GlitchData : VitalGlitchDataType;
	variable  PPCS0PLBRDDBUS54_GlitchData : VitalGlitchDataType;
	variable  PPCS0PLBRDDBUS55_GlitchData : VitalGlitchDataType;
	variable  PPCS0PLBRDDBUS56_GlitchData : VitalGlitchDataType;
	variable  PPCS0PLBRDDBUS57_GlitchData : VitalGlitchDataType;
	variable  PPCS0PLBRDDBUS58_GlitchData : VitalGlitchDataType;
	variable  PPCS0PLBRDDBUS59_GlitchData : VitalGlitchDataType;
	variable  PPCS0PLBRDDBUS60_GlitchData : VitalGlitchDataType;
	variable  PPCS0PLBRDDBUS61_GlitchData : VitalGlitchDataType;
	variable  PPCS0PLBRDDBUS62_GlitchData : VitalGlitchDataType;
	variable  PPCS0PLBRDDBUS63_GlitchData : VitalGlitchDataType;
	variable  PPCS0PLBRDDBUS64_GlitchData : VitalGlitchDataType;
	variable  PPCS0PLBRDDBUS65_GlitchData : VitalGlitchDataType;
	variable  PPCS0PLBRDDBUS66_GlitchData : VitalGlitchDataType;
	variable  PPCS0PLBRDDBUS67_GlitchData : VitalGlitchDataType;
	variable  PPCS0PLBRDDBUS68_GlitchData : VitalGlitchDataType;
	variable  PPCS0PLBRDDBUS69_GlitchData : VitalGlitchDataType;
	variable  PPCS0PLBRDDBUS70_GlitchData : VitalGlitchDataType;
	variable  PPCS0PLBRDDBUS71_GlitchData : VitalGlitchDataType;
	variable  PPCS0PLBRDDBUS72_GlitchData : VitalGlitchDataType;
	variable  PPCS0PLBRDDBUS73_GlitchData : VitalGlitchDataType;
	variable  PPCS0PLBRDDBUS74_GlitchData : VitalGlitchDataType;
	variable  PPCS0PLBRDDBUS75_GlitchData : VitalGlitchDataType;
	variable  PPCS0PLBRDDBUS76_GlitchData : VitalGlitchDataType;
	variable  PPCS0PLBRDDBUS77_GlitchData : VitalGlitchDataType;
	variable  PPCS0PLBRDDBUS78_GlitchData : VitalGlitchDataType;
	variable  PPCS0PLBRDDBUS79_GlitchData : VitalGlitchDataType;
	variable  PPCS0PLBRDDBUS80_GlitchData : VitalGlitchDataType;
	variable  PPCS0PLBRDDBUS81_GlitchData : VitalGlitchDataType;
	variable  PPCS0PLBRDDBUS82_GlitchData : VitalGlitchDataType;
	variable  PPCS0PLBRDDBUS83_GlitchData : VitalGlitchDataType;
	variable  PPCS0PLBRDDBUS84_GlitchData : VitalGlitchDataType;
	variable  PPCS0PLBRDDBUS85_GlitchData : VitalGlitchDataType;
	variable  PPCS0PLBRDDBUS86_GlitchData : VitalGlitchDataType;
	variable  PPCS0PLBRDDBUS87_GlitchData : VitalGlitchDataType;
	variable  PPCS0PLBRDDBUS88_GlitchData : VitalGlitchDataType;
	variable  PPCS0PLBRDDBUS89_GlitchData : VitalGlitchDataType;
	variable  PPCS0PLBRDDBUS90_GlitchData : VitalGlitchDataType;
	variable  PPCS0PLBRDDBUS91_GlitchData : VitalGlitchDataType;
	variable  PPCS0PLBRDDBUS92_GlitchData : VitalGlitchDataType;
	variable  PPCS0PLBRDDBUS93_GlitchData : VitalGlitchDataType;
	variable  PPCS0PLBRDDBUS94_GlitchData : VitalGlitchDataType;
	variable  PPCS0PLBRDDBUS95_GlitchData : VitalGlitchDataType;
	variable  PPCS0PLBRDDBUS96_GlitchData : VitalGlitchDataType;
	variable  PPCS0PLBRDDBUS97_GlitchData : VitalGlitchDataType;
	variable  PPCS0PLBRDDBUS98_GlitchData : VitalGlitchDataType;
	variable  PPCS0PLBRDDBUS99_GlitchData : VitalGlitchDataType;
	variable  PPCS0PLBRDDBUS100_GlitchData : VitalGlitchDataType;
	variable  PPCS0PLBRDDBUS101_GlitchData : VitalGlitchDataType;
	variable  PPCS0PLBRDDBUS102_GlitchData : VitalGlitchDataType;
	variable  PPCS0PLBRDDBUS103_GlitchData : VitalGlitchDataType;
	variable  PPCS0PLBRDDBUS104_GlitchData : VitalGlitchDataType;
	variable  PPCS0PLBRDDBUS105_GlitchData : VitalGlitchDataType;
	variable  PPCS0PLBRDDBUS106_GlitchData : VitalGlitchDataType;
	variable  PPCS0PLBRDDBUS107_GlitchData : VitalGlitchDataType;
	variable  PPCS0PLBRDDBUS108_GlitchData : VitalGlitchDataType;
	variable  PPCS0PLBRDDBUS109_GlitchData : VitalGlitchDataType;
	variable  PPCS0PLBRDDBUS110_GlitchData : VitalGlitchDataType;
	variable  PPCS0PLBRDDBUS111_GlitchData : VitalGlitchDataType;
	variable  PPCS0PLBRDDBUS112_GlitchData : VitalGlitchDataType;
	variable  PPCS0PLBRDDBUS113_GlitchData : VitalGlitchDataType;
	variable  PPCS0PLBRDDBUS114_GlitchData : VitalGlitchDataType;
	variable  PPCS0PLBRDDBUS115_GlitchData : VitalGlitchDataType;
	variable  PPCS0PLBRDDBUS116_GlitchData : VitalGlitchDataType;
	variable  PPCS0PLBRDDBUS117_GlitchData : VitalGlitchDataType;
	variable  PPCS0PLBRDDBUS118_GlitchData : VitalGlitchDataType;
	variable  PPCS0PLBRDDBUS119_GlitchData : VitalGlitchDataType;
	variable  PPCS0PLBRDDBUS120_GlitchData : VitalGlitchDataType;
	variable  PPCS0PLBRDDBUS121_GlitchData : VitalGlitchDataType;
	variable  PPCS0PLBRDDBUS122_GlitchData : VitalGlitchDataType;
	variable  PPCS0PLBRDDBUS123_GlitchData : VitalGlitchDataType;
	variable  PPCS0PLBRDDBUS124_GlitchData : VitalGlitchDataType;
	variable  PPCS0PLBRDDBUS125_GlitchData : VitalGlitchDataType;
	variable  PPCS0PLBRDDBUS126_GlitchData : VitalGlitchDataType;
	variable  PPCS0PLBRDDBUS127_GlitchData : VitalGlitchDataType;
	variable  PPCS0PLBRDWDADDR0_GlitchData : VitalGlitchDataType;
	variable  PPCS0PLBRDWDADDR1_GlitchData : VitalGlitchDataType;
	variable  PPCS0PLBRDWDADDR2_GlitchData : VitalGlitchDataType;
	variable  PPCS0PLBRDWDADDR3_GlitchData : VitalGlitchDataType;
	variable  PPCS0PLBREARBITRATE_GlitchData : VitalGlitchDataType;
	variable  PPCS0PLBSSIZE0_GlitchData : VitalGlitchDataType;
	variable  PPCS0PLBSSIZE1_GlitchData : VitalGlitchDataType;
	variable  PPCS0PLBWAIT_GlitchData : VitalGlitchDataType;
	variable  PPCS0PLBWRBTERM_GlitchData : VitalGlitchDataType;
	variable  PPCS0PLBWRCOMP_GlitchData : VitalGlitchDataType;
	variable  PPCS0PLBWRDACK_GlitchData : VitalGlitchDataType;
	variable  PPCS1PLBADDRACK_GlitchData : VitalGlitchDataType;
	variable  PPCS1PLBMBUSY0_GlitchData : VitalGlitchDataType;
	variable  PPCS1PLBMBUSY1_GlitchData : VitalGlitchDataType;
	variable  PPCS1PLBMBUSY2_GlitchData : VitalGlitchDataType;
	variable  PPCS1PLBMBUSY3_GlitchData : VitalGlitchDataType;
	variable  PPCS1PLBMIRQ0_GlitchData : VitalGlitchDataType;
	variable  PPCS1PLBMIRQ1_GlitchData : VitalGlitchDataType;
	variable  PPCS1PLBMIRQ2_GlitchData : VitalGlitchDataType;
	variable  PPCS1PLBMIRQ3_GlitchData : VitalGlitchDataType;
	variable  PPCS1PLBMRDERR0_GlitchData : VitalGlitchDataType;
	variable  PPCS1PLBMRDERR1_GlitchData : VitalGlitchDataType;
	variable  PPCS1PLBMRDERR2_GlitchData : VitalGlitchDataType;
	variable  PPCS1PLBMRDERR3_GlitchData : VitalGlitchDataType;
	variable  PPCS1PLBMWRERR0_GlitchData : VitalGlitchDataType;
	variable  PPCS1PLBMWRERR1_GlitchData : VitalGlitchDataType;
	variable  PPCS1PLBMWRERR2_GlitchData : VitalGlitchDataType;
	variable  PPCS1PLBMWRERR3_GlitchData : VitalGlitchDataType;
	variable  PPCS1PLBRDBTERM_GlitchData : VitalGlitchDataType;
	variable  PPCS1PLBRDCOMP_GlitchData : VitalGlitchDataType;
	variable  PPCS1PLBRDDACK_GlitchData : VitalGlitchDataType;
	variable  PPCS1PLBRDDBUS0_GlitchData : VitalGlitchDataType;
	variable  PPCS1PLBRDDBUS1_GlitchData : VitalGlitchDataType;
	variable  PPCS1PLBRDDBUS2_GlitchData : VitalGlitchDataType;
	variable  PPCS1PLBRDDBUS3_GlitchData : VitalGlitchDataType;
	variable  PPCS1PLBRDDBUS4_GlitchData : VitalGlitchDataType;
	variable  PPCS1PLBRDDBUS5_GlitchData : VitalGlitchDataType;
	variable  PPCS1PLBRDDBUS6_GlitchData : VitalGlitchDataType;
	variable  PPCS1PLBRDDBUS7_GlitchData : VitalGlitchDataType;
	variable  PPCS1PLBRDDBUS8_GlitchData : VitalGlitchDataType;
	variable  PPCS1PLBRDDBUS9_GlitchData : VitalGlitchDataType;
	variable  PPCS1PLBRDDBUS10_GlitchData : VitalGlitchDataType;
	variable  PPCS1PLBRDDBUS11_GlitchData : VitalGlitchDataType;
	variable  PPCS1PLBRDDBUS12_GlitchData : VitalGlitchDataType;
	variable  PPCS1PLBRDDBUS13_GlitchData : VitalGlitchDataType;
	variable  PPCS1PLBRDDBUS14_GlitchData : VitalGlitchDataType;
	variable  PPCS1PLBRDDBUS15_GlitchData : VitalGlitchDataType;
	variable  PPCS1PLBRDDBUS16_GlitchData : VitalGlitchDataType;
	variable  PPCS1PLBRDDBUS17_GlitchData : VitalGlitchDataType;
	variable  PPCS1PLBRDDBUS18_GlitchData : VitalGlitchDataType;
	variable  PPCS1PLBRDDBUS19_GlitchData : VitalGlitchDataType;
	variable  PPCS1PLBRDDBUS20_GlitchData : VitalGlitchDataType;
	variable  PPCS1PLBRDDBUS21_GlitchData : VitalGlitchDataType;
	variable  PPCS1PLBRDDBUS22_GlitchData : VitalGlitchDataType;
	variable  PPCS1PLBRDDBUS23_GlitchData : VitalGlitchDataType;
	variable  PPCS1PLBRDDBUS24_GlitchData : VitalGlitchDataType;
	variable  PPCS1PLBRDDBUS25_GlitchData : VitalGlitchDataType;
	variable  PPCS1PLBRDDBUS26_GlitchData : VitalGlitchDataType;
	variable  PPCS1PLBRDDBUS27_GlitchData : VitalGlitchDataType;
	variable  PPCS1PLBRDDBUS28_GlitchData : VitalGlitchDataType;
	variable  PPCS1PLBRDDBUS29_GlitchData : VitalGlitchDataType;
	variable  PPCS1PLBRDDBUS30_GlitchData : VitalGlitchDataType;
	variable  PPCS1PLBRDDBUS31_GlitchData : VitalGlitchDataType;
	variable  PPCS1PLBRDDBUS32_GlitchData : VitalGlitchDataType;
	variable  PPCS1PLBRDDBUS33_GlitchData : VitalGlitchDataType;
	variable  PPCS1PLBRDDBUS34_GlitchData : VitalGlitchDataType;
	variable  PPCS1PLBRDDBUS35_GlitchData : VitalGlitchDataType;
	variable  PPCS1PLBRDDBUS36_GlitchData : VitalGlitchDataType;
	variable  PPCS1PLBRDDBUS37_GlitchData : VitalGlitchDataType;
	variable  PPCS1PLBRDDBUS38_GlitchData : VitalGlitchDataType;
	variable  PPCS1PLBRDDBUS39_GlitchData : VitalGlitchDataType;
	variable  PPCS1PLBRDDBUS40_GlitchData : VitalGlitchDataType;
	variable  PPCS1PLBRDDBUS41_GlitchData : VitalGlitchDataType;
	variable  PPCS1PLBRDDBUS42_GlitchData : VitalGlitchDataType;
	variable  PPCS1PLBRDDBUS43_GlitchData : VitalGlitchDataType;
	variable  PPCS1PLBRDDBUS44_GlitchData : VitalGlitchDataType;
	variable  PPCS1PLBRDDBUS45_GlitchData : VitalGlitchDataType;
	variable  PPCS1PLBRDDBUS46_GlitchData : VitalGlitchDataType;
	variable  PPCS1PLBRDDBUS47_GlitchData : VitalGlitchDataType;
	variable  PPCS1PLBRDDBUS48_GlitchData : VitalGlitchDataType;
	variable  PPCS1PLBRDDBUS49_GlitchData : VitalGlitchDataType;
	variable  PPCS1PLBRDDBUS50_GlitchData : VitalGlitchDataType;
	variable  PPCS1PLBRDDBUS51_GlitchData : VitalGlitchDataType;
	variable  PPCS1PLBRDDBUS52_GlitchData : VitalGlitchDataType;
	variable  PPCS1PLBRDDBUS53_GlitchData : VitalGlitchDataType;
	variable  PPCS1PLBRDDBUS54_GlitchData : VitalGlitchDataType;
	variable  PPCS1PLBRDDBUS55_GlitchData : VitalGlitchDataType;
	variable  PPCS1PLBRDDBUS56_GlitchData : VitalGlitchDataType;
	variable  PPCS1PLBRDDBUS57_GlitchData : VitalGlitchDataType;
	variable  PPCS1PLBRDDBUS58_GlitchData : VitalGlitchDataType;
	variable  PPCS1PLBRDDBUS59_GlitchData : VitalGlitchDataType;
	variable  PPCS1PLBRDDBUS60_GlitchData : VitalGlitchDataType;
	variable  PPCS1PLBRDDBUS61_GlitchData : VitalGlitchDataType;
	variable  PPCS1PLBRDDBUS62_GlitchData : VitalGlitchDataType;
	variable  PPCS1PLBRDDBUS63_GlitchData : VitalGlitchDataType;
	variable  PPCS1PLBRDDBUS64_GlitchData : VitalGlitchDataType;
	variable  PPCS1PLBRDDBUS65_GlitchData : VitalGlitchDataType;
	variable  PPCS1PLBRDDBUS66_GlitchData : VitalGlitchDataType;
	variable  PPCS1PLBRDDBUS67_GlitchData : VitalGlitchDataType;
	variable  PPCS1PLBRDDBUS68_GlitchData : VitalGlitchDataType;
	variable  PPCS1PLBRDDBUS69_GlitchData : VitalGlitchDataType;
	variable  PPCS1PLBRDDBUS70_GlitchData : VitalGlitchDataType;
	variable  PPCS1PLBRDDBUS71_GlitchData : VitalGlitchDataType;
	variable  PPCS1PLBRDDBUS72_GlitchData : VitalGlitchDataType;
	variable  PPCS1PLBRDDBUS73_GlitchData : VitalGlitchDataType;
	variable  PPCS1PLBRDDBUS74_GlitchData : VitalGlitchDataType;
	variable  PPCS1PLBRDDBUS75_GlitchData : VitalGlitchDataType;
	variable  PPCS1PLBRDDBUS76_GlitchData : VitalGlitchDataType;
	variable  PPCS1PLBRDDBUS77_GlitchData : VitalGlitchDataType;
	variable  PPCS1PLBRDDBUS78_GlitchData : VitalGlitchDataType;
	variable  PPCS1PLBRDDBUS79_GlitchData : VitalGlitchDataType;
	variable  PPCS1PLBRDDBUS80_GlitchData : VitalGlitchDataType;
	variable  PPCS1PLBRDDBUS81_GlitchData : VitalGlitchDataType;
	variable  PPCS1PLBRDDBUS82_GlitchData : VitalGlitchDataType;
	variable  PPCS1PLBRDDBUS83_GlitchData : VitalGlitchDataType;
	variable  PPCS1PLBRDDBUS84_GlitchData : VitalGlitchDataType;
	variable  PPCS1PLBRDDBUS85_GlitchData : VitalGlitchDataType;
	variable  PPCS1PLBRDDBUS86_GlitchData : VitalGlitchDataType;
	variable  PPCS1PLBRDDBUS87_GlitchData : VitalGlitchDataType;
	variable  PPCS1PLBRDDBUS88_GlitchData : VitalGlitchDataType;
	variable  PPCS1PLBRDDBUS89_GlitchData : VitalGlitchDataType;
	variable  PPCS1PLBRDDBUS90_GlitchData : VitalGlitchDataType;
	variable  PPCS1PLBRDDBUS91_GlitchData : VitalGlitchDataType;
	variable  PPCS1PLBRDDBUS92_GlitchData : VitalGlitchDataType;
	variable  PPCS1PLBRDDBUS93_GlitchData : VitalGlitchDataType;
	variable  PPCS1PLBRDDBUS94_GlitchData : VitalGlitchDataType;
	variable  PPCS1PLBRDDBUS95_GlitchData : VitalGlitchDataType;
	variable  PPCS1PLBRDDBUS96_GlitchData : VitalGlitchDataType;
	variable  PPCS1PLBRDDBUS97_GlitchData : VitalGlitchDataType;
	variable  PPCS1PLBRDDBUS98_GlitchData : VitalGlitchDataType;
	variable  PPCS1PLBRDDBUS99_GlitchData : VitalGlitchDataType;
	variable  PPCS1PLBRDDBUS100_GlitchData : VitalGlitchDataType;
	variable  PPCS1PLBRDDBUS101_GlitchData : VitalGlitchDataType;
	variable  PPCS1PLBRDDBUS102_GlitchData : VitalGlitchDataType;
	variable  PPCS1PLBRDDBUS103_GlitchData : VitalGlitchDataType;
	variable  PPCS1PLBRDDBUS104_GlitchData : VitalGlitchDataType;
	variable  PPCS1PLBRDDBUS105_GlitchData : VitalGlitchDataType;
	variable  PPCS1PLBRDDBUS106_GlitchData : VitalGlitchDataType;
	variable  PPCS1PLBRDDBUS107_GlitchData : VitalGlitchDataType;
	variable  PPCS1PLBRDDBUS108_GlitchData : VitalGlitchDataType;
	variable  PPCS1PLBRDDBUS109_GlitchData : VitalGlitchDataType;
	variable  PPCS1PLBRDDBUS110_GlitchData : VitalGlitchDataType;
	variable  PPCS1PLBRDDBUS111_GlitchData : VitalGlitchDataType;
	variable  PPCS1PLBRDDBUS112_GlitchData : VitalGlitchDataType;
	variable  PPCS1PLBRDDBUS113_GlitchData : VitalGlitchDataType;
	variable  PPCS1PLBRDDBUS114_GlitchData : VitalGlitchDataType;
	variable  PPCS1PLBRDDBUS115_GlitchData : VitalGlitchDataType;
	variable  PPCS1PLBRDDBUS116_GlitchData : VitalGlitchDataType;
	variable  PPCS1PLBRDDBUS117_GlitchData : VitalGlitchDataType;
	variable  PPCS1PLBRDDBUS118_GlitchData : VitalGlitchDataType;
	variable  PPCS1PLBRDDBUS119_GlitchData : VitalGlitchDataType;
	variable  PPCS1PLBRDDBUS120_GlitchData : VitalGlitchDataType;
	variable  PPCS1PLBRDDBUS121_GlitchData : VitalGlitchDataType;
	variable  PPCS1PLBRDDBUS122_GlitchData : VitalGlitchDataType;
	variable  PPCS1PLBRDDBUS123_GlitchData : VitalGlitchDataType;
	variable  PPCS1PLBRDDBUS124_GlitchData : VitalGlitchDataType;
	variable  PPCS1PLBRDDBUS125_GlitchData : VitalGlitchDataType;
	variable  PPCS1PLBRDDBUS126_GlitchData : VitalGlitchDataType;
	variable  PPCS1PLBRDDBUS127_GlitchData : VitalGlitchDataType;
	variable  PPCS1PLBRDWDADDR0_GlitchData : VitalGlitchDataType;
	variable  PPCS1PLBRDWDADDR1_GlitchData : VitalGlitchDataType;
	variable  PPCS1PLBRDWDADDR2_GlitchData : VitalGlitchDataType;
	variable  PPCS1PLBRDWDADDR3_GlitchData : VitalGlitchDataType;
	variable  PPCS1PLBREARBITRATE_GlitchData : VitalGlitchDataType;
	variable  PPCS1PLBSSIZE0_GlitchData : VitalGlitchDataType;
	variable  PPCS1PLBSSIZE1_GlitchData : VitalGlitchDataType;
	variable  PPCS1PLBWAIT_GlitchData : VitalGlitchDataType;
	variable  PPCS1PLBWRBTERM_GlitchData : VitalGlitchDataType;
	variable  PPCS1PLBWRCOMP_GlitchData : VitalGlitchDataType;
	variable  PPCS1PLBWRDACK_GlitchData : VitalGlitchDataType;
	variable  APUFCMDECFPUOP_GlitchData : VitalGlitchDataType;
	variable  APUFCMDECLDSTXFERSIZE0_GlitchData : VitalGlitchDataType;
	variable  APUFCMDECLDSTXFERSIZE1_GlitchData : VitalGlitchDataType;
	variable  APUFCMDECLDSTXFERSIZE2_GlitchData : VitalGlitchDataType;
	variable  APUFCMDECLOAD_GlitchData : VitalGlitchDataType;
	variable  APUFCMDECNONAUTON_GlitchData : VitalGlitchDataType;
	variable  APUFCMDECSTORE_GlitchData : VitalGlitchDataType;
	variable  APUFCMDECUDI0_GlitchData : VitalGlitchDataType;
	variable  APUFCMDECUDI1_GlitchData : VitalGlitchDataType;
	variable  APUFCMDECUDI2_GlitchData : VitalGlitchDataType;
	variable  APUFCMDECUDI3_GlitchData : VitalGlitchDataType;
	variable  APUFCMDECUDIVALID_GlitchData : VitalGlitchDataType;
	variable  APUFCMENDIAN_GlitchData : VitalGlitchDataType;
	variable  APUFCMFLUSH_GlitchData : VitalGlitchDataType;
	variable  APUFCMINSTRUCTION0_GlitchData : VitalGlitchDataType;
	variable  APUFCMINSTRUCTION1_GlitchData : VitalGlitchDataType;
	variable  APUFCMINSTRUCTION2_GlitchData : VitalGlitchDataType;
	variable  APUFCMINSTRUCTION3_GlitchData : VitalGlitchDataType;
	variable  APUFCMINSTRUCTION4_GlitchData : VitalGlitchDataType;
	variable  APUFCMINSTRUCTION5_GlitchData : VitalGlitchDataType;
	variable  APUFCMINSTRUCTION6_GlitchData : VitalGlitchDataType;
	variable  APUFCMINSTRUCTION7_GlitchData : VitalGlitchDataType;
	variable  APUFCMINSTRUCTION8_GlitchData : VitalGlitchDataType;
	variable  APUFCMINSTRUCTION9_GlitchData : VitalGlitchDataType;
	variable  APUFCMINSTRUCTION10_GlitchData : VitalGlitchDataType;
	variable  APUFCMINSTRUCTION11_GlitchData : VitalGlitchDataType;
	variable  APUFCMINSTRUCTION12_GlitchData : VitalGlitchDataType;
	variable  APUFCMINSTRUCTION13_GlitchData : VitalGlitchDataType;
	variable  APUFCMINSTRUCTION14_GlitchData : VitalGlitchDataType;
	variable  APUFCMINSTRUCTION15_GlitchData : VitalGlitchDataType;
	variable  APUFCMINSTRUCTION16_GlitchData : VitalGlitchDataType;
	variable  APUFCMINSTRUCTION17_GlitchData : VitalGlitchDataType;
	variable  APUFCMINSTRUCTION18_GlitchData : VitalGlitchDataType;
	variable  APUFCMINSTRUCTION19_GlitchData : VitalGlitchDataType;
	variable  APUFCMINSTRUCTION20_GlitchData : VitalGlitchDataType;
	variable  APUFCMINSTRUCTION21_GlitchData : VitalGlitchDataType;
	variable  APUFCMINSTRUCTION22_GlitchData : VitalGlitchDataType;
	variable  APUFCMINSTRUCTION23_GlitchData : VitalGlitchDataType;
	variable  APUFCMINSTRUCTION24_GlitchData : VitalGlitchDataType;
	variable  APUFCMINSTRUCTION25_GlitchData : VitalGlitchDataType;
	variable  APUFCMINSTRUCTION26_GlitchData : VitalGlitchDataType;
	variable  APUFCMINSTRUCTION27_GlitchData : VitalGlitchDataType;
	variable  APUFCMINSTRUCTION28_GlitchData : VitalGlitchDataType;
	variable  APUFCMINSTRUCTION29_GlitchData : VitalGlitchDataType;
	variable  APUFCMINSTRUCTION30_GlitchData : VitalGlitchDataType;
	variable  APUFCMINSTRUCTION31_GlitchData : VitalGlitchDataType;
	variable  APUFCMINSTRVALID_GlitchData : VitalGlitchDataType;
	variable  APUFCMLOADBYTEADDR0_GlitchData : VitalGlitchDataType;
	variable  APUFCMLOADBYTEADDR1_GlitchData : VitalGlitchDataType;
	variable  APUFCMLOADBYTEADDR2_GlitchData : VitalGlitchDataType;
	variable  APUFCMLOADBYTEADDR3_GlitchData : VitalGlitchDataType;
	variable  APUFCMLOADDATA0_GlitchData : VitalGlitchDataType;
	variable  APUFCMLOADDATA1_GlitchData : VitalGlitchDataType;
	variable  APUFCMLOADDATA2_GlitchData : VitalGlitchDataType;
	variable  APUFCMLOADDATA3_GlitchData : VitalGlitchDataType;
	variable  APUFCMLOADDATA4_GlitchData : VitalGlitchDataType;
	variable  APUFCMLOADDATA5_GlitchData : VitalGlitchDataType;
	variable  APUFCMLOADDATA6_GlitchData : VitalGlitchDataType;
	variable  APUFCMLOADDATA7_GlitchData : VitalGlitchDataType;
	variable  APUFCMLOADDATA8_GlitchData : VitalGlitchDataType;
	variable  APUFCMLOADDATA9_GlitchData : VitalGlitchDataType;
	variable  APUFCMLOADDATA10_GlitchData : VitalGlitchDataType;
	variable  APUFCMLOADDATA11_GlitchData : VitalGlitchDataType;
	variable  APUFCMLOADDATA12_GlitchData : VitalGlitchDataType;
	variable  APUFCMLOADDATA13_GlitchData : VitalGlitchDataType;
	variable  APUFCMLOADDATA14_GlitchData : VitalGlitchDataType;
	variable  APUFCMLOADDATA15_GlitchData : VitalGlitchDataType;
	variable  APUFCMLOADDATA16_GlitchData : VitalGlitchDataType;
	variable  APUFCMLOADDATA17_GlitchData : VitalGlitchDataType;
	variable  APUFCMLOADDATA18_GlitchData : VitalGlitchDataType;
	variable  APUFCMLOADDATA19_GlitchData : VitalGlitchDataType;
	variable  APUFCMLOADDATA20_GlitchData : VitalGlitchDataType;
	variable  APUFCMLOADDATA21_GlitchData : VitalGlitchDataType;
	variable  APUFCMLOADDATA22_GlitchData : VitalGlitchDataType;
	variable  APUFCMLOADDATA23_GlitchData : VitalGlitchDataType;
	variable  APUFCMLOADDATA24_GlitchData : VitalGlitchDataType;
	variable  APUFCMLOADDATA25_GlitchData : VitalGlitchDataType;
	variable  APUFCMLOADDATA26_GlitchData : VitalGlitchDataType;
	variable  APUFCMLOADDATA27_GlitchData : VitalGlitchDataType;
	variable  APUFCMLOADDATA28_GlitchData : VitalGlitchDataType;
	variable  APUFCMLOADDATA29_GlitchData : VitalGlitchDataType;
	variable  APUFCMLOADDATA30_GlitchData : VitalGlitchDataType;
	variable  APUFCMLOADDATA31_GlitchData : VitalGlitchDataType;
	variable  APUFCMLOADDATA32_GlitchData : VitalGlitchDataType;
	variable  APUFCMLOADDATA33_GlitchData : VitalGlitchDataType;
	variable  APUFCMLOADDATA34_GlitchData : VitalGlitchDataType;
	variable  APUFCMLOADDATA35_GlitchData : VitalGlitchDataType;
	variable  APUFCMLOADDATA36_GlitchData : VitalGlitchDataType;
	variable  APUFCMLOADDATA37_GlitchData : VitalGlitchDataType;
	variable  APUFCMLOADDATA38_GlitchData : VitalGlitchDataType;
	variable  APUFCMLOADDATA39_GlitchData : VitalGlitchDataType;
	variable  APUFCMLOADDATA40_GlitchData : VitalGlitchDataType;
	variable  APUFCMLOADDATA41_GlitchData : VitalGlitchDataType;
	variable  APUFCMLOADDATA42_GlitchData : VitalGlitchDataType;
	variable  APUFCMLOADDATA43_GlitchData : VitalGlitchDataType;
	variable  APUFCMLOADDATA44_GlitchData : VitalGlitchDataType;
	variable  APUFCMLOADDATA45_GlitchData : VitalGlitchDataType;
	variable  APUFCMLOADDATA46_GlitchData : VitalGlitchDataType;
	variable  APUFCMLOADDATA47_GlitchData : VitalGlitchDataType;
	variable  APUFCMLOADDATA48_GlitchData : VitalGlitchDataType;
	variable  APUFCMLOADDATA49_GlitchData : VitalGlitchDataType;
	variable  APUFCMLOADDATA50_GlitchData : VitalGlitchDataType;
	variable  APUFCMLOADDATA51_GlitchData : VitalGlitchDataType;
	variable  APUFCMLOADDATA52_GlitchData : VitalGlitchDataType;
	variable  APUFCMLOADDATA53_GlitchData : VitalGlitchDataType;
	variable  APUFCMLOADDATA54_GlitchData : VitalGlitchDataType;
	variable  APUFCMLOADDATA55_GlitchData : VitalGlitchDataType;
	variable  APUFCMLOADDATA56_GlitchData : VitalGlitchDataType;
	variable  APUFCMLOADDATA57_GlitchData : VitalGlitchDataType;
	variable  APUFCMLOADDATA58_GlitchData : VitalGlitchDataType;
	variable  APUFCMLOADDATA59_GlitchData : VitalGlitchDataType;
	variable  APUFCMLOADDATA60_GlitchData : VitalGlitchDataType;
	variable  APUFCMLOADDATA61_GlitchData : VitalGlitchDataType;
	variable  APUFCMLOADDATA62_GlitchData : VitalGlitchDataType;
	variable  APUFCMLOADDATA63_GlitchData : VitalGlitchDataType;
	variable  APUFCMLOADDATA64_GlitchData : VitalGlitchDataType;
	variable  APUFCMLOADDATA65_GlitchData : VitalGlitchDataType;
	variable  APUFCMLOADDATA66_GlitchData : VitalGlitchDataType;
	variable  APUFCMLOADDATA67_GlitchData : VitalGlitchDataType;
	variable  APUFCMLOADDATA68_GlitchData : VitalGlitchDataType;
	variable  APUFCMLOADDATA69_GlitchData : VitalGlitchDataType;
	variable  APUFCMLOADDATA70_GlitchData : VitalGlitchDataType;
	variable  APUFCMLOADDATA71_GlitchData : VitalGlitchDataType;
	variable  APUFCMLOADDATA72_GlitchData : VitalGlitchDataType;
	variable  APUFCMLOADDATA73_GlitchData : VitalGlitchDataType;
	variable  APUFCMLOADDATA74_GlitchData : VitalGlitchDataType;
	variable  APUFCMLOADDATA75_GlitchData : VitalGlitchDataType;
	variable  APUFCMLOADDATA76_GlitchData : VitalGlitchDataType;
	variable  APUFCMLOADDATA77_GlitchData : VitalGlitchDataType;
	variable  APUFCMLOADDATA78_GlitchData : VitalGlitchDataType;
	variable  APUFCMLOADDATA79_GlitchData : VitalGlitchDataType;
	variable  APUFCMLOADDATA80_GlitchData : VitalGlitchDataType;
	variable  APUFCMLOADDATA81_GlitchData : VitalGlitchDataType;
	variable  APUFCMLOADDATA82_GlitchData : VitalGlitchDataType;
	variable  APUFCMLOADDATA83_GlitchData : VitalGlitchDataType;
	variable  APUFCMLOADDATA84_GlitchData : VitalGlitchDataType;
	variable  APUFCMLOADDATA85_GlitchData : VitalGlitchDataType;
	variable  APUFCMLOADDATA86_GlitchData : VitalGlitchDataType;
	variable  APUFCMLOADDATA87_GlitchData : VitalGlitchDataType;
	variable  APUFCMLOADDATA88_GlitchData : VitalGlitchDataType;
	variable  APUFCMLOADDATA89_GlitchData : VitalGlitchDataType;
	variable  APUFCMLOADDATA90_GlitchData : VitalGlitchDataType;
	variable  APUFCMLOADDATA91_GlitchData : VitalGlitchDataType;
	variable  APUFCMLOADDATA92_GlitchData : VitalGlitchDataType;
	variable  APUFCMLOADDATA93_GlitchData : VitalGlitchDataType;
	variable  APUFCMLOADDATA94_GlitchData : VitalGlitchDataType;
	variable  APUFCMLOADDATA95_GlitchData : VitalGlitchDataType;
	variable  APUFCMLOADDATA96_GlitchData : VitalGlitchDataType;
	variable  APUFCMLOADDATA97_GlitchData : VitalGlitchDataType;
	variable  APUFCMLOADDATA98_GlitchData : VitalGlitchDataType;
	variable  APUFCMLOADDATA99_GlitchData : VitalGlitchDataType;
	variable  APUFCMLOADDATA100_GlitchData : VitalGlitchDataType;
	variable  APUFCMLOADDATA101_GlitchData : VitalGlitchDataType;
	variable  APUFCMLOADDATA102_GlitchData : VitalGlitchDataType;
	variable  APUFCMLOADDATA103_GlitchData : VitalGlitchDataType;
	variable  APUFCMLOADDATA104_GlitchData : VitalGlitchDataType;
	variable  APUFCMLOADDATA105_GlitchData : VitalGlitchDataType;
	variable  APUFCMLOADDATA106_GlitchData : VitalGlitchDataType;
	variable  APUFCMLOADDATA107_GlitchData : VitalGlitchDataType;
	variable  APUFCMLOADDATA108_GlitchData : VitalGlitchDataType;
	variable  APUFCMLOADDATA109_GlitchData : VitalGlitchDataType;
	variable  APUFCMLOADDATA110_GlitchData : VitalGlitchDataType;
	variable  APUFCMLOADDATA111_GlitchData : VitalGlitchDataType;
	variable  APUFCMLOADDATA112_GlitchData : VitalGlitchDataType;
	variable  APUFCMLOADDATA113_GlitchData : VitalGlitchDataType;
	variable  APUFCMLOADDATA114_GlitchData : VitalGlitchDataType;
	variable  APUFCMLOADDATA115_GlitchData : VitalGlitchDataType;
	variable  APUFCMLOADDATA116_GlitchData : VitalGlitchDataType;
	variable  APUFCMLOADDATA117_GlitchData : VitalGlitchDataType;
	variable  APUFCMLOADDATA118_GlitchData : VitalGlitchDataType;
	variable  APUFCMLOADDATA119_GlitchData : VitalGlitchDataType;
	variable  APUFCMLOADDATA120_GlitchData : VitalGlitchDataType;
	variable  APUFCMLOADDATA121_GlitchData : VitalGlitchDataType;
	variable  APUFCMLOADDATA122_GlitchData : VitalGlitchDataType;
	variable  APUFCMLOADDATA123_GlitchData : VitalGlitchDataType;
	variable  APUFCMLOADDATA124_GlitchData : VitalGlitchDataType;
	variable  APUFCMLOADDATA125_GlitchData : VitalGlitchDataType;
	variable  APUFCMLOADDATA126_GlitchData : VitalGlitchDataType;
	variable  APUFCMLOADDATA127_GlitchData : VitalGlitchDataType;
	variable  APUFCMLOADDVALID_GlitchData : VitalGlitchDataType;
	variable  APUFCMMSRFE0_GlitchData : VitalGlitchDataType;
	variable  APUFCMMSRFE1_GlitchData : VitalGlitchDataType;
	variable  APUFCMNEXTINSTRREADY_GlitchData : VitalGlitchDataType;
	variable  APUFCMOPERANDVALID_GlitchData : VitalGlitchDataType;
	variable  APUFCMRADATA0_GlitchData : VitalGlitchDataType;
	variable  APUFCMRADATA1_GlitchData : VitalGlitchDataType;
	variable  APUFCMRADATA2_GlitchData : VitalGlitchDataType;
	variable  APUFCMRADATA3_GlitchData : VitalGlitchDataType;
	variable  APUFCMRADATA4_GlitchData : VitalGlitchDataType;
	variable  APUFCMRADATA5_GlitchData : VitalGlitchDataType;
	variable  APUFCMRADATA6_GlitchData : VitalGlitchDataType;
	variable  APUFCMRADATA7_GlitchData : VitalGlitchDataType;
	variable  APUFCMRADATA8_GlitchData : VitalGlitchDataType;
	variable  APUFCMRADATA9_GlitchData : VitalGlitchDataType;
	variable  APUFCMRADATA10_GlitchData : VitalGlitchDataType;
	variable  APUFCMRADATA11_GlitchData : VitalGlitchDataType;
	variable  APUFCMRADATA12_GlitchData : VitalGlitchDataType;
	variable  APUFCMRADATA13_GlitchData : VitalGlitchDataType;
	variable  APUFCMRADATA14_GlitchData : VitalGlitchDataType;
	variable  APUFCMRADATA15_GlitchData : VitalGlitchDataType;
	variable  APUFCMRADATA16_GlitchData : VitalGlitchDataType;
	variable  APUFCMRADATA17_GlitchData : VitalGlitchDataType;
	variable  APUFCMRADATA18_GlitchData : VitalGlitchDataType;
	variable  APUFCMRADATA19_GlitchData : VitalGlitchDataType;
	variable  APUFCMRADATA20_GlitchData : VitalGlitchDataType;
	variable  APUFCMRADATA21_GlitchData : VitalGlitchDataType;
	variable  APUFCMRADATA22_GlitchData : VitalGlitchDataType;
	variable  APUFCMRADATA23_GlitchData : VitalGlitchDataType;
	variable  APUFCMRADATA24_GlitchData : VitalGlitchDataType;
	variable  APUFCMRADATA25_GlitchData : VitalGlitchDataType;
	variable  APUFCMRADATA26_GlitchData : VitalGlitchDataType;
	variable  APUFCMRADATA27_GlitchData : VitalGlitchDataType;
	variable  APUFCMRADATA28_GlitchData : VitalGlitchDataType;
	variable  APUFCMRADATA29_GlitchData : VitalGlitchDataType;
	variable  APUFCMRADATA30_GlitchData : VitalGlitchDataType;
	variable  APUFCMRADATA31_GlitchData : VitalGlitchDataType;
	variable  APUFCMRBDATA0_GlitchData : VitalGlitchDataType;
	variable  APUFCMRBDATA1_GlitchData : VitalGlitchDataType;
	variable  APUFCMRBDATA2_GlitchData : VitalGlitchDataType;
	variable  APUFCMRBDATA3_GlitchData : VitalGlitchDataType;
	variable  APUFCMRBDATA4_GlitchData : VitalGlitchDataType;
	variable  APUFCMRBDATA5_GlitchData : VitalGlitchDataType;
	variable  APUFCMRBDATA6_GlitchData : VitalGlitchDataType;
	variable  APUFCMRBDATA7_GlitchData : VitalGlitchDataType;
	variable  APUFCMRBDATA8_GlitchData : VitalGlitchDataType;
	variable  APUFCMRBDATA9_GlitchData : VitalGlitchDataType;
	variable  APUFCMRBDATA10_GlitchData : VitalGlitchDataType;
	variable  APUFCMRBDATA11_GlitchData : VitalGlitchDataType;
	variable  APUFCMRBDATA12_GlitchData : VitalGlitchDataType;
	variable  APUFCMRBDATA13_GlitchData : VitalGlitchDataType;
	variable  APUFCMRBDATA14_GlitchData : VitalGlitchDataType;
	variable  APUFCMRBDATA15_GlitchData : VitalGlitchDataType;
	variable  APUFCMRBDATA16_GlitchData : VitalGlitchDataType;
	variable  APUFCMRBDATA17_GlitchData : VitalGlitchDataType;
	variable  APUFCMRBDATA18_GlitchData : VitalGlitchDataType;
	variable  APUFCMRBDATA19_GlitchData : VitalGlitchDataType;
	variable  APUFCMRBDATA20_GlitchData : VitalGlitchDataType;
	variable  APUFCMRBDATA21_GlitchData : VitalGlitchDataType;
	variable  APUFCMRBDATA22_GlitchData : VitalGlitchDataType;
	variable  APUFCMRBDATA23_GlitchData : VitalGlitchDataType;
	variable  APUFCMRBDATA24_GlitchData : VitalGlitchDataType;
	variable  APUFCMRBDATA25_GlitchData : VitalGlitchDataType;
	variable  APUFCMRBDATA26_GlitchData : VitalGlitchDataType;
	variable  APUFCMRBDATA27_GlitchData : VitalGlitchDataType;
	variable  APUFCMRBDATA28_GlitchData : VitalGlitchDataType;
	variable  APUFCMRBDATA29_GlitchData : VitalGlitchDataType;
	variable  APUFCMRBDATA30_GlitchData : VitalGlitchDataType;
	variable  APUFCMRBDATA31_GlitchData : VitalGlitchDataType;
	variable  APUFCMWRITEBACKOK_GlitchData : VitalGlitchDataType;
	variable  C440CPMCORESLEEPREQ_GlitchData : VitalGlitchDataType;
	variable  C440CPMDECIRPTREQ_GlitchData : VitalGlitchDataType;
	variable  C440CPMFITIRPTREQ_GlitchData : VitalGlitchDataType;
	variable  C440CPMMSRCE_GlitchData : VitalGlitchDataType;
	variable  C440CPMMSREE_GlitchData : VitalGlitchDataType;
	variable  C440CPMTIMERRESETREQ_GlitchData : VitalGlitchDataType;
	variable  C440CPMWDIRPTREQ_GlitchData : VitalGlitchDataType;
	variable  C440DBGSYSTEMCONTROL0_GlitchData : VitalGlitchDataType;
	variable  C440DBGSYSTEMCONTROL1_GlitchData : VitalGlitchDataType;
	variable  C440DBGSYSTEMCONTROL2_GlitchData : VitalGlitchDataType;
	variable  C440DBGSYSTEMCONTROL3_GlitchData : VitalGlitchDataType;
	variable  C440DBGSYSTEMCONTROL4_GlitchData : VitalGlitchDataType;
	variable  C440DBGSYSTEMCONTROL5_GlitchData : VitalGlitchDataType;
	variable  C440DBGSYSTEMCONTROL6_GlitchData : VitalGlitchDataType;
	variable  C440DBGSYSTEMCONTROL7_GlitchData : VitalGlitchDataType;
	variable  C440JTGTDO_GlitchData : VitalGlitchDataType;
	variable  C440JTGTDOEN_GlitchData : VitalGlitchDataType;
	variable  C440MACHINECHECK_GlitchData : VitalGlitchDataType;
	variable  C440RSTCHIPRESETREQ_GlitchData : VitalGlitchDataType;
	variable  C440RSTCORERESETREQ_GlitchData : VitalGlitchDataType;
	variable  C440RSTSYSTEMRESETREQ_GlitchData : VitalGlitchDataType;
	variable  C440TRCBRANCHSTATUS0_GlitchData : VitalGlitchDataType;
	variable  C440TRCBRANCHSTATUS1_GlitchData : VitalGlitchDataType;
	variable  C440TRCBRANCHSTATUS2_GlitchData : VitalGlitchDataType;
	variable  C440TRCCYCLE_GlitchData : VitalGlitchDataType;
	variable  C440TRCEXECUTIONSTATUS0_GlitchData : VitalGlitchDataType;
	variable  C440TRCEXECUTIONSTATUS1_GlitchData : VitalGlitchDataType;
	variable  C440TRCEXECUTIONSTATUS2_GlitchData : VitalGlitchDataType;
	variable  C440TRCEXECUTIONSTATUS3_GlitchData : VitalGlitchDataType;
	variable  C440TRCEXECUTIONSTATUS4_GlitchData : VitalGlitchDataType;
	variable  C440TRCTRACESTATUS0_GlitchData : VitalGlitchDataType;
	variable  C440TRCTRACESTATUS1_GlitchData : VitalGlitchDataType;
	variable  C440TRCTRACESTATUS2_GlitchData : VitalGlitchDataType;
	variable  C440TRCTRACESTATUS3_GlitchData : VitalGlitchDataType;
	variable  C440TRCTRACESTATUS4_GlitchData : VitalGlitchDataType;
	variable  C440TRCTRACESTATUS5_GlitchData : VitalGlitchDataType;
	variable  C440TRCTRACESTATUS6_GlitchData : VitalGlitchDataType;
	variable  C440TRCTRIGGEREVENTOUT_GlitchData : VitalGlitchDataType;
	variable  C440TRCTRIGGEREVENTTYPE0_GlitchData : VitalGlitchDataType;
	variable  C440TRCTRIGGEREVENTTYPE1_GlitchData : VitalGlitchDataType;
	variable  C440TRCTRIGGEREVENTTYPE2_GlitchData : VitalGlitchDataType;
	variable  C440TRCTRIGGEREVENTTYPE3_GlitchData : VitalGlitchDataType;
	variable  C440TRCTRIGGEREVENTTYPE4_GlitchData : VitalGlitchDataType;
	variable  C440TRCTRIGGEREVENTTYPE5_GlitchData : VitalGlitchDataType;
	variable  C440TRCTRIGGEREVENTTYPE6_GlitchData : VitalGlitchDataType;
	variable  C440TRCTRIGGEREVENTTYPE7_GlitchData : VitalGlitchDataType;
	variable  C440TRCTRIGGEREVENTTYPE8_GlitchData : VitalGlitchDataType;
	variable  C440TRCTRIGGEREVENTTYPE9_GlitchData : VitalGlitchDataType;
	variable  C440TRCTRIGGEREVENTTYPE10_GlitchData : VitalGlitchDataType;
	variable  C440TRCTRIGGEREVENTTYPE11_GlitchData : VitalGlitchDataType;
	variable  C440TRCTRIGGEREVENTTYPE12_GlitchData : VitalGlitchDataType;
	variable  C440TRCTRIGGEREVENTTYPE13_GlitchData : VitalGlitchDataType;
	variable  MIMCADDRESS0_GlitchData : VitalGlitchDataType;
	variable  MIMCADDRESS1_GlitchData : VitalGlitchDataType;
	variable  MIMCADDRESS2_GlitchData : VitalGlitchDataType;
	variable  MIMCADDRESS3_GlitchData : VitalGlitchDataType;
	variable  MIMCADDRESS4_GlitchData : VitalGlitchDataType;
	variable  MIMCADDRESS5_GlitchData : VitalGlitchDataType;
	variable  MIMCADDRESS6_GlitchData : VitalGlitchDataType;
	variable  MIMCADDRESS7_GlitchData : VitalGlitchDataType;
	variable  MIMCADDRESS8_GlitchData : VitalGlitchDataType;
	variable  MIMCADDRESS9_GlitchData : VitalGlitchDataType;
	variable  MIMCADDRESS10_GlitchData : VitalGlitchDataType;
	variable  MIMCADDRESS11_GlitchData : VitalGlitchDataType;
	variable  MIMCADDRESS12_GlitchData : VitalGlitchDataType;
	variable  MIMCADDRESS13_GlitchData : VitalGlitchDataType;
	variable  MIMCADDRESS14_GlitchData : VitalGlitchDataType;
	variable  MIMCADDRESS15_GlitchData : VitalGlitchDataType;
	variable  MIMCADDRESS16_GlitchData : VitalGlitchDataType;
	variable  MIMCADDRESS17_GlitchData : VitalGlitchDataType;
	variable  MIMCADDRESS18_GlitchData : VitalGlitchDataType;
	variable  MIMCADDRESS19_GlitchData : VitalGlitchDataType;
	variable  MIMCADDRESS20_GlitchData : VitalGlitchDataType;
	variable  MIMCADDRESS21_GlitchData : VitalGlitchDataType;
	variable  MIMCADDRESS22_GlitchData : VitalGlitchDataType;
	variable  MIMCADDRESS23_GlitchData : VitalGlitchDataType;
	variable  MIMCADDRESS24_GlitchData : VitalGlitchDataType;
	variable  MIMCADDRESS25_GlitchData : VitalGlitchDataType;
	variable  MIMCADDRESS26_GlitchData : VitalGlitchDataType;
	variable  MIMCADDRESS27_GlitchData : VitalGlitchDataType;
	variable  MIMCADDRESS28_GlitchData : VitalGlitchDataType;
	variable  MIMCADDRESS29_GlitchData : VitalGlitchDataType;
	variable  MIMCADDRESS30_GlitchData : VitalGlitchDataType;
	variable  MIMCADDRESS31_GlitchData : VitalGlitchDataType;
	variable  MIMCADDRESS32_GlitchData : VitalGlitchDataType;
	variable  MIMCADDRESS33_GlitchData : VitalGlitchDataType;
	variable  MIMCADDRESS34_GlitchData : VitalGlitchDataType;
	variable  MIMCADDRESS35_GlitchData : VitalGlitchDataType;
	variable  MIMCADDRESSVALID_GlitchData : VitalGlitchDataType;
	variable  MIMCBANKCONFLICT_GlitchData : VitalGlitchDataType;
	variable  MIMCBYTEENABLE0_GlitchData : VitalGlitchDataType;
	variable  MIMCBYTEENABLE1_GlitchData : VitalGlitchDataType;
	variable  MIMCBYTEENABLE2_GlitchData : VitalGlitchDataType;
	variable  MIMCBYTEENABLE3_GlitchData : VitalGlitchDataType;
	variable  MIMCBYTEENABLE4_GlitchData : VitalGlitchDataType;
	variable  MIMCBYTEENABLE5_GlitchData : VitalGlitchDataType;
	variable  MIMCBYTEENABLE6_GlitchData : VitalGlitchDataType;
	variable  MIMCBYTEENABLE7_GlitchData : VitalGlitchDataType;
	variable  MIMCBYTEENABLE8_GlitchData : VitalGlitchDataType;
	variable  MIMCBYTEENABLE9_GlitchData : VitalGlitchDataType;
	variable  MIMCBYTEENABLE10_GlitchData : VitalGlitchDataType;
	variable  MIMCBYTEENABLE11_GlitchData : VitalGlitchDataType;
	variable  MIMCBYTEENABLE12_GlitchData : VitalGlitchDataType;
	variable  MIMCBYTEENABLE13_GlitchData : VitalGlitchDataType;
	variable  MIMCBYTEENABLE14_GlitchData : VitalGlitchDataType;
	variable  MIMCBYTEENABLE15_GlitchData : VitalGlitchDataType;
	variable  MIMCREADNOTWRITE_GlitchData : VitalGlitchDataType;
	variable  MIMCROWCONFLICT_GlitchData : VitalGlitchDataType;
	variable  MIMCWRITEDATA0_GlitchData : VitalGlitchDataType;
	variable  MIMCWRITEDATA1_GlitchData : VitalGlitchDataType;
	variable  MIMCWRITEDATA2_GlitchData : VitalGlitchDataType;
	variable  MIMCWRITEDATA3_GlitchData : VitalGlitchDataType;
	variable  MIMCWRITEDATA4_GlitchData : VitalGlitchDataType;
	variable  MIMCWRITEDATA5_GlitchData : VitalGlitchDataType;
	variable  MIMCWRITEDATA6_GlitchData : VitalGlitchDataType;
	variable  MIMCWRITEDATA7_GlitchData : VitalGlitchDataType;
	variable  MIMCWRITEDATA8_GlitchData : VitalGlitchDataType;
	variable  MIMCWRITEDATA9_GlitchData : VitalGlitchDataType;
	variable  MIMCWRITEDATA10_GlitchData : VitalGlitchDataType;
	variable  MIMCWRITEDATA11_GlitchData : VitalGlitchDataType;
	variable  MIMCWRITEDATA12_GlitchData : VitalGlitchDataType;
	variable  MIMCWRITEDATA13_GlitchData : VitalGlitchDataType;
	variable  MIMCWRITEDATA14_GlitchData : VitalGlitchDataType;
	variable  MIMCWRITEDATA15_GlitchData : VitalGlitchDataType;
	variable  MIMCWRITEDATA16_GlitchData : VitalGlitchDataType;
	variable  MIMCWRITEDATA17_GlitchData : VitalGlitchDataType;
	variable  MIMCWRITEDATA18_GlitchData : VitalGlitchDataType;
	variable  MIMCWRITEDATA19_GlitchData : VitalGlitchDataType;
	variable  MIMCWRITEDATA20_GlitchData : VitalGlitchDataType;
	variable  MIMCWRITEDATA21_GlitchData : VitalGlitchDataType;
	variable  MIMCWRITEDATA22_GlitchData : VitalGlitchDataType;
	variable  MIMCWRITEDATA23_GlitchData : VitalGlitchDataType;
	variable  MIMCWRITEDATA24_GlitchData : VitalGlitchDataType;
	variable  MIMCWRITEDATA25_GlitchData : VitalGlitchDataType;
	variable  MIMCWRITEDATA26_GlitchData : VitalGlitchDataType;
	variable  MIMCWRITEDATA27_GlitchData : VitalGlitchDataType;
	variable  MIMCWRITEDATA28_GlitchData : VitalGlitchDataType;
	variable  MIMCWRITEDATA29_GlitchData : VitalGlitchDataType;
	variable  MIMCWRITEDATA30_GlitchData : VitalGlitchDataType;
	variable  MIMCWRITEDATA31_GlitchData : VitalGlitchDataType;
	variable  MIMCWRITEDATA32_GlitchData : VitalGlitchDataType;
	variable  MIMCWRITEDATA33_GlitchData : VitalGlitchDataType;
	variable  MIMCWRITEDATA34_GlitchData : VitalGlitchDataType;
	variable  MIMCWRITEDATA35_GlitchData : VitalGlitchDataType;
	variable  MIMCWRITEDATA36_GlitchData : VitalGlitchDataType;
	variable  MIMCWRITEDATA37_GlitchData : VitalGlitchDataType;
	variable  MIMCWRITEDATA38_GlitchData : VitalGlitchDataType;
	variable  MIMCWRITEDATA39_GlitchData : VitalGlitchDataType;
	variable  MIMCWRITEDATA40_GlitchData : VitalGlitchDataType;
	variable  MIMCWRITEDATA41_GlitchData : VitalGlitchDataType;
	variable  MIMCWRITEDATA42_GlitchData : VitalGlitchDataType;
	variable  MIMCWRITEDATA43_GlitchData : VitalGlitchDataType;
	variable  MIMCWRITEDATA44_GlitchData : VitalGlitchDataType;
	variable  MIMCWRITEDATA45_GlitchData : VitalGlitchDataType;
	variable  MIMCWRITEDATA46_GlitchData : VitalGlitchDataType;
	variable  MIMCWRITEDATA47_GlitchData : VitalGlitchDataType;
	variable  MIMCWRITEDATA48_GlitchData : VitalGlitchDataType;
	variable  MIMCWRITEDATA49_GlitchData : VitalGlitchDataType;
	variable  MIMCWRITEDATA50_GlitchData : VitalGlitchDataType;
	variable  MIMCWRITEDATA51_GlitchData : VitalGlitchDataType;
	variable  MIMCWRITEDATA52_GlitchData : VitalGlitchDataType;
	variable  MIMCWRITEDATA53_GlitchData : VitalGlitchDataType;
	variable  MIMCWRITEDATA54_GlitchData : VitalGlitchDataType;
	variable  MIMCWRITEDATA55_GlitchData : VitalGlitchDataType;
	variable  MIMCWRITEDATA56_GlitchData : VitalGlitchDataType;
	variable  MIMCWRITEDATA57_GlitchData : VitalGlitchDataType;
	variable  MIMCWRITEDATA58_GlitchData : VitalGlitchDataType;
	variable  MIMCWRITEDATA59_GlitchData : VitalGlitchDataType;
	variable  MIMCWRITEDATA60_GlitchData : VitalGlitchDataType;
	variable  MIMCWRITEDATA61_GlitchData : VitalGlitchDataType;
	variable  MIMCWRITEDATA62_GlitchData : VitalGlitchDataType;
	variable  MIMCWRITEDATA63_GlitchData : VitalGlitchDataType;
	variable  MIMCWRITEDATA64_GlitchData : VitalGlitchDataType;
	variable  MIMCWRITEDATA65_GlitchData : VitalGlitchDataType;
	variable  MIMCWRITEDATA66_GlitchData : VitalGlitchDataType;
	variable  MIMCWRITEDATA67_GlitchData : VitalGlitchDataType;
	variable  MIMCWRITEDATA68_GlitchData : VitalGlitchDataType;
	variable  MIMCWRITEDATA69_GlitchData : VitalGlitchDataType;
	variable  MIMCWRITEDATA70_GlitchData : VitalGlitchDataType;
	variable  MIMCWRITEDATA71_GlitchData : VitalGlitchDataType;
	variable  MIMCWRITEDATA72_GlitchData : VitalGlitchDataType;
	variable  MIMCWRITEDATA73_GlitchData : VitalGlitchDataType;
	variable  MIMCWRITEDATA74_GlitchData : VitalGlitchDataType;
	variable  MIMCWRITEDATA75_GlitchData : VitalGlitchDataType;
	variable  MIMCWRITEDATA76_GlitchData : VitalGlitchDataType;
	variable  MIMCWRITEDATA77_GlitchData : VitalGlitchDataType;
	variable  MIMCWRITEDATA78_GlitchData : VitalGlitchDataType;
	variable  MIMCWRITEDATA79_GlitchData : VitalGlitchDataType;
	variable  MIMCWRITEDATA80_GlitchData : VitalGlitchDataType;
	variable  MIMCWRITEDATA81_GlitchData : VitalGlitchDataType;
	variable  MIMCWRITEDATA82_GlitchData : VitalGlitchDataType;
	variable  MIMCWRITEDATA83_GlitchData : VitalGlitchDataType;
	variable  MIMCWRITEDATA84_GlitchData : VitalGlitchDataType;
	variable  MIMCWRITEDATA85_GlitchData : VitalGlitchDataType;
	variable  MIMCWRITEDATA86_GlitchData : VitalGlitchDataType;
	variable  MIMCWRITEDATA87_GlitchData : VitalGlitchDataType;
	variable  MIMCWRITEDATA88_GlitchData : VitalGlitchDataType;
	variable  MIMCWRITEDATA89_GlitchData : VitalGlitchDataType;
	variable  MIMCWRITEDATA90_GlitchData : VitalGlitchDataType;
	variable  MIMCWRITEDATA91_GlitchData : VitalGlitchDataType;
	variable  MIMCWRITEDATA92_GlitchData : VitalGlitchDataType;
	variable  MIMCWRITEDATA93_GlitchData : VitalGlitchDataType;
	variable  MIMCWRITEDATA94_GlitchData : VitalGlitchDataType;
	variable  MIMCWRITEDATA95_GlitchData : VitalGlitchDataType;
	variable  MIMCWRITEDATA96_GlitchData : VitalGlitchDataType;
	variable  MIMCWRITEDATA97_GlitchData : VitalGlitchDataType;
	variable  MIMCWRITEDATA98_GlitchData : VitalGlitchDataType;
	variable  MIMCWRITEDATA99_GlitchData : VitalGlitchDataType;
	variable  MIMCWRITEDATA100_GlitchData : VitalGlitchDataType;
	variable  MIMCWRITEDATA101_GlitchData : VitalGlitchDataType;
	variable  MIMCWRITEDATA102_GlitchData : VitalGlitchDataType;
	variable  MIMCWRITEDATA103_GlitchData : VitalGlitchDataType;
	variable  MIMCWRITEDATA104_GlitchData : VitalGlitchDataType;
	variable  MIMCWRITEDATA105_GlitchData : VitalGlitchDataType;
	variable  MIMCWRITEDATA106_GlitchData : VitalGlitchDataType;
	variable  MIMCWRITEDATA107_GlitchData : VitalGlitchDataType;
	variable  MIMCWRITEDATA108_GlitchData : VitalGlitchDataType;
	variable  MIMCWRITEDATA109_GlitchData : VitalGlitchDataType;
	variable  MIMCWRITEDATA110_GlitchData : VitalGlitchDataType;
	variable  MIMCWRITEDATA111_GlitchData : VitalGlitchDataType;
	variable  MIMCWRITEDATA112_GlitchData : VitalGlitchDataType;
	variable  MIMCWRITEDATA113_GlitchData : VitalGlitchDataType;
	variable  MIMCWRITEDATA114_GlitchData : VitalGlitchDataType;
	variable  MIMCWRITEDATA115_GlitchData : VitalGlitchDataType;
	variable  MIMCWRITEDATA116_GlitchData : VitalGlitchDataType;
	variable  MIMCWRITEDATA117_GlitchData : VitalGlitchDataType;
	variable  MIMCWRITEDATA118_GlitchData : VitalGlitchDataType;
	variable  MIMCWRITEDATA119_GlitchData : VitalGlitchDataType;
	variable  MIMCWRITEDATA120_GlitchData : VitalGlitchDataType;
	variable  MIMCWRITEDATA121_GlitchData : VitalGlitchDataType;
	variable  MIMCWRITEDATA122_GlitchData : VitalGlitchDataType;
	variable  MIMCWRITEDATA123_GlitchData : VitalGlitchDataType;
	variable  MIMCWRITEDATA124_GlitchData : VitalGlitchDataType;
	variable  MIMCWRITEDATA125_GlitchData : VitalGlitchDataType;
	variable  MIMCWRITEDATA126_GlitchData : VitalGlitchDataType;
	variable  MIMCWRITEDATA127_GlitchData : VitalGlitchDataType;
	variable  MIMCWRITEDATAVALID_GlitchData : VitalGlitchDataType;
	variable  PPCCPMINTERCONNECTBUSY_GlitchData : VitalGlitchDataType;
	variable  PPCDSDCRACK_GlitchData : VitalGlitchDataType;
	variable  PPCDSDCRTIMEOUTWAIT_GlitchData : VitalGlitchDataType;
	variable  PPCDSDCRDBUSIN0_GlitchData : VitalGlitchDataType;
	variable  PPCDSDCRDBUSIN1_GlitchData : VitalGlitchDataType;
	variable  PPCDSDCRDBUSIN2_GlitchData : VitalGlitchDataType;
	variable  PPCDSDCRDBUSIN3_GlitchData : VitalGlitchDataType;
	variable  PPCDSDCRDBUSIN4_GlitchData : VitalGlitchDataType;
	variable  PPCDSDCRDBUSIN5_GlitchData : VitalGlitchDataType;
	variable  PPCDSDCRDBUSIN6_GlitchData : VitalGlitchDataType;
	variable  PPCDSDCRDBUSIN7_GlitchData : VitalGlitchDataType;
	variable  PPCDSDCRDBUSIN8_GlitchData : VitalGlitchDataType;
	variable  PPCDSDCRDBUSIN9_GlitchData : VitalGlitchDataType;
	variable  PPCDSDCRDBUSIN10_GlitchData : VitalGlitchDataType;
	variable  PPCDSDCRDBUSIN11_GlitchData : VitalGlitchDataType;
	variable  PPCDSDCRDBUSIN12_GlitchData : VitalGlitchDataType;
	variable  PPCDSDCRDBUSIN13_GlitchData : VitalGlitchDataType;
	variable  PPCDSDCRDBUSIN14_GlitchData : VitalGlitchDataType;
	variable  PPCDSDCRDBUSIN15_GlitchData : VitalGlitchDataType;
	variable  PPCDSDCRDBUSIN16_GlitchData : VitalGlitchDataType;
	variable  PPCDSDCRDBUSIN17_GlitchData : VitalGlitchDataType;
	variable  PPCDSDCRDBUSIN18_GlitchData : VitalGlitchDataType;
	variable  PPCDSDCRDBUSIN19_GlitchData : VitalGlitchDataType;
	variable  PPCDSDCRDBUSIN20_GlitchData : VitalGlitchDataType;
	variable  PPCDSDCRDBUSIN21_GlitchData : VitalGlitchDataType;
	variable  PPCDSDCRDBUSIN22_GlitchData : VitalGlitchDataType;
	variable  PPCDSDCRDBUSIN23_GlitchData : VitalGlitchDataType;
	variable  PPCDSDCRDBUSIN24_GlitchData : VitalGlitchDataType;
	variable  PPCDSDCRDBUSIN25_GlitchData : VitalGlitchDataType;
	variable  PPCDSDCRDBUSIN26_GlitchData : VitalGlitchDataType;
	variable  PPCDSDCRDBUSIN27_GlitchData : VitalGlitchDataType;
	variable  PPCDSDCRDBUSIN28_GlitchData : VitalGlitchDataType;
	variable  PPCDSDCRDBUSIN29_GlitchData : VitalGlitchDataType;
	variable  PPCDSDCRDBUSIN30_GlitchData : VitalGlitchDataType;
	variable  PPCDSDCRDBUSIN31_GlitchData : VitalGlitchDataType;
	variable  PPCEICINTERCONNECTIRQ_GlitchData : VitalGlitchDataType;
begin

	VitalPathDelay01
	(
	OutSignal     => DMA0LLRSTENGINEACK,
	GlitchData    => DMA0LLRSTENGINEACK_GlitchData,
	OutSignalName => "DMA0LLRSTENGINEACK",
	OutTemp       => DMA0LLRSTENGINEACK_OUT,
	Paths         => (0 => (CPMDMA0LLCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => DMA0LLRXDSTRDYN,
	GlitchData    => DMA0LLRXDSTRDYN_GlitchData,
	OutSignalName => "DMA0LLRXDSTRDYN",
	OutTemp       => DMA0LLRXDSTRDYN_OUT,
	Paths         => (0 => (CPMDMA0LLCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => DMA0LLTXD(0),
	GlitchData    => DMA0LLTXD0_GlitchData,
	OutSignalName => "DMA0LLTXD(0)",
	OutTemp       => DMA0LLTXD_OUT(0),
	Paths         => (0 => (CPMDMA0LLCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => DMA0LLTXD(1),
	GlitchData    => DMA0LLTXD1_GlitchData,
	OutSignalName => "DMA0LLTXD(1)",
	OutTemp       => DMA0LLTXD_OUT(1),
	Paths         => (0 => (CPMDMA0LLCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => DMA0LLTXD(2),
	GlitchData    => DMA0LLTXD2_GlitchData,
	OutSignalName => "DMA0LLTXD(2)",
	OutTemp       => DMA0LLTXD_OUT(2),
	Paths         => (0 => (CPMDMA0LLCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => DMA0LLTXD(3),
	GlitchData    => DMA0LLTXD3_GlitchData,
	OutSignalName => "DMA0LLTXD(3)",
	OutTemp       => DMA0LLTXD_OUT(3),
	Paths         => (0 => (CPMDMA0LLCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => DMA0LLTXD(4),
	GlitchData    => DMA0LLTXD4_GlitchData,
	OutSignalName => "DMA0LLTXD(4)",
	OutTemp       => DMA0LLTXD_OUT(4),
	Paths         => (0 => (CPMDMA0LLCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => DMA0LLTXD(5),
	GlitchData    => DMA0LLTXD5_GlitchData,
	OutSignalName => "DMA0LLTXD(5)",
	OutTemp       => DMA0LLTXD_OUT(5),
	Paths         => (0 => (CPMDMA0LLCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => DMA0LLTXD(6),
	GlitchData    => DMA0LLTXD6_GlitchData,
	OutSignalName => "DMA0LLTXD(6)",
	OutTemp       => DMA0LLTXD_OUT(6),
	Paths         => (0 => (CPMDMA0LLCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => DMA0LLTXD(7),
	GlitchData    => DMA0LLTXD7_GlitchData,
	OutSignalName => "DMA0LLTXD(7)",
	OutTemp       => DMA0LLTXD_OUT(7),
	Paths         => (0 => (CPMDMA0LLCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => DMA0LLTXD(8),
	GlitchData    => DMA0LLTXD8_GlitchData,
	OutSignalName => "DMA0LLTXD(8)",
	OutTemp       => DMA0LLTXD_OUT(8),
	Paths         => (0 => (CPMDMA0LLCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => DMA0LLTXD(9),
	GlitchData    => DMA0LLTXD9_GlitchData,
	OutSignalName => "DMA0LLTXD(9)",
	OutTemp       => DMA0LLTXD_OUT(9),
	Paths         => (0 => (CPMDMA0LLCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => DMA0LLTXD(10),
	GlitchData    => DMA0LLTXD10_GlitchData,
	OutSignalName => "DMA0LLTXD(10)",
	OutTemp       => DMA0LLTXD_OUT(10),
	Paths         => (0 => (CPMDMA0LLCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => DMA0LLTXD(11),
	GlitchData    => DMA0LLTXD11_GlitchData,
	OutSignalName => "DMA0LLTXD(11)",
	OutTemp       => DMA0LLTXD_OUT(11),
	Paths         => (0 => (CPMDMA0LLCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => DMA0LLTXD(12),
	GlitchData    => DMA0LLTXD12_GlitchData,
	OutSignalName => "DMA0LLTXD(12)",
	OutTemp       => DMA0LLTXD_OUT(12),
	Paths         => (0 => (CPMDMA0LLCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => DMA0LLTXD(13),
	GlitchData    => DMA0LLTXD13_GlitchData,
	OutSignalName => "DMA0LLTXD(13)",
	OutTemp       => DMA0LLTXD_OUT(13),
	Paths         => (0 => (CPMDMA0LLCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => DMA0LLTXD(14),
	GlitchData    => DMA0LLTXD14_GlitchData,
	OutSignalName => "DMA0LLTXD(14)",
	OutTemp       => DMA0LLTXD_OUT(14),
	Paths         => (0 => (CPMDMA0LLCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => DMA0LLTXD(15),
	GlitchData    => DMA0LLTXD15_GlitchData,
	OutSignalName => "DMA0LLTXD(15)",
	OutTemp       => DMA0LLTXD_OUT(15),
	Paths         => (0 => (CPMDMA0LLCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => DMA0LLTXD(16),
	GlitchData    => DMA0LLTXD16_GlitchData,
	OutSignalName => "DMA0LLTXD(16)",
	OutTemp       => DMA0LLTXD_OUT(16),
	Paths         => (0 => (CPMDMA0LLCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => DMA0LLTXD(17),
	GlitchData    => DMA0LLTXD17_GlitchData,
	OutSignalName => "DMA0LLTXD(17)",
	OutTemp       => DMA0LLTXD_OUT(17),
	Paths         => (0 => (CPMDMA0LLCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => DMA0LLTXD(18),
	GlitchData    => DMA0LLTXD18_GlitchData,
	OutSignalName => "DMA0LLTXD(18)",
	OutTemp       => DMA0LLTXD_OUT(18),
	Paths         => (0 => (CPMDMA0LLCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => DMA0LLTXD(19),
	GlitchData    => DMA0LLTXD19_GlitchData,
	OutSignalName => "DMA0LLTXD(19)",
	OutTemp       => DMA0LLTXD_OUT(19),
	Paths         => (0 => (CPMDMA0LLCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => DMA0LLTXD(20),
	GlitchData    => DMA0LLTXD20_GlitchData,
	OutSignalName => "DMA0LLTXD(20)",
	OutTemp       => DMA0LLTXD_OUT(20),
	Paths         => (0 => (CPMDMA0LLCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => DMA0LLTXD(21),
	GlitchData    => DMA0LLTXD21_GlitchData,
	OutSignalName => "DMA0LLTXD(21)",
	OutTemp       => DMA0LLTXD_OUT(21),
	Paths         => (0 => (CPMDMA0LLCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => DMA0LLTXD(22),
	GlitchData    => DMA0LLTXD22_GlitchData,
	OutSignalName => "DMA0LLTXD(22)",
	OutTemp       => DMA0LLTXD_OUT(22),
	Paths         => (0 => (CPMDMA0LLCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => DMA0LLTXD(23),
	GlitchData    => DMA0LLTXD23_GlitchData,
	OutSignalName => "DMA0LLTXD(23)",
	OutTemp       => DMA0LLTXD_OUT(23),
	Paths         => (0 => (CPMDMA0LLCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => DMA0LLTXD(24),
	GlitchData    => DMA0LLTXD24_GlitchData,
	OutSignalName => "DMA0LLTXD(24)",
	OutTemp       => DMA0LLTXD_OUT(24),
	Paths         => (0 => (CPMDMA0LLCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => DMA0LLTXD(25),
	GlitchData    => DMA0LLTXD25_GlitchData,
	OutSignalName => "DMA0LLTXD(25)",
	OutTemp       => DMA0LLTXD_OUT(25),
	Paths         => (0 => (CPMDMA0LLCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => DMA0LLTXD(26),
	GlitchData    => DMA0LLTXD26_GlitchData,
	OutSignalName => "DMA0LLTXD(26)",
	OutTemp       => DMA0LLTXD_OUT(26),
	Paths         => (0 => (CPMDMA0LLCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => DMA0LLTXD(27),
	GlitchData    => DMA0LLTXD27_GlitchData,
	OutSignalName => "DMA0LLTXD(27)",
	OutTemp       => DMA0LLTXD_OUT(27),
	Paths         => (0 => (CPMDMA0LLCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => DMA0LLTXD(28),
	GlitchData    => DMA0LLTXD28_GlitchData,
	OutSignalName => "DMA0LLTXD(28)",
	OutTemp       => DMA0LLTXD_OUT(28),
	Paths         => (0 => (CPMDMA0LLCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => DMA0LLTXD(29),
	GlitchData    => DMA0LLTXD29_GlitchData,
	OutSignalName => "DMA0LLTXD(29)",
	OutTemp       => DMA0LLTXD_OUT(29),
	Paths         => (0 => (CPMDMA0LLCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => DMA0LLTXD(30),
	GlitchData    => DMA0LLTXD30_GlitchData,
	OutSignalName => "DMA0LLTXD(30)",
	OutTemp       => DMA0LLTXD_OUT(30),
	Paths         => (0 => (CPMDMA0LLCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => DMA0LLTXD(31),
	GlitchData    => DMA0LLTXD31_GlitchData,
	OutSignalName => "DMA0LLTXD(31)",
	OutTemp       => DMA0LLTXD_OUT(31),
	Paths         => (0 => (CPMDMA0LLCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => DMA0LLTXEOFN,
	GlitchData    => DMA0LLTXEOFN_GlitchData,
	OutSignalName => "DMA0LLTXEOFN",
	OutTemp       => DMA0LLTXEOFN_OUT,
	Paths         => (0 => (CPMDMA0LLCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => DMA0LLTXEOPN,
	GlitchData    => DMA0LLTXEOPN_GlitchData,
	OutSignalName => "DMA0LLTXEOPN",
	OutTemp       => DMA0LLTXEOPN_OUT,
	Paths         => (0 => (CPMDMA0LLCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => DMA0LLTXREM(0),
	GlitchData    => DMA0LLTXREM0_GlitchData,
	OutSignalName => "DMA0LLTXREM(0)",
	OutTemp       => DMA0LLTXREM_OUT(0),
	Paths         => (0 => (CPMDMA0LLCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => DMA0LLTXREM(1),
	GlitchData    => DMA0LLTXREM1_GlitchData,
	OutSignalName => "DMA0LLTXREM(1)",
	OutTemp       => DMA0LLTXREM_OUT(1),
	Paths         => (0 => (CPMDMA0LLCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => DMA0LLTXREM(2),
	GlitchData    => DMA0LLTXREM2_GlitchData,
	OutSignalName => "DMA0LLTXREM(2)",
	OutTemp       => DMA0LLTXREM_OUT(2),
	Paths         => (0 => (CPMDMA0LLCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => DMA0LLTXREM(3),
	GlitchData    => DMA0LLTXREM3_GlitchData,
	OutSignalName => "DMA0LLTXREM(3)",
	OutTemp       => DMA0LLTXREM_OUT(3),
	Paths         => (0 => (CPMDMA0LLCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => DMA0LLTXSOFN,
	GlitchData    => DMA0LLTXSOFN_GlitchData,
	OutSignalName => "DMA0LLTXSOFN",
	OutTemp       => DMA0LLTXSOFN_OUT,
	Paths         => (0 => (CPMDMA0LLCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => DMA0LLTXSOPN,
	GlitchData    => DMA0LLTXSOPN_GlitchData,
	OutSignalName => "DMA0LLTXSOPN",
	OutTemp       => DMA0LLTXSOPN_OUT,
	Paths         => (0 => (CPMDMA0LLCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => DMA0LLTXSRCRDYN,
	GlitchData    => DMA0LLTXSRCRDYN_GlitchData,
	OutSignalName => "DMA0LLTXSRCRDYN",
	OutTemp       => DMA0LLTXSRCRDYN_OUT,
	Paths         => (0 => (CPMDMA0LLCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => DMA0RXIRQ,
	GlitchData    => DMA0RXIRQ_GlitchData,
	OutSignalName => "DMA0RXIRQ",
	OutTemp       => DMA0RXIRQ_OUT,
	Paths         => (0 => (CPMDMA0LLCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => DMA0TXIRQ,
	GlitchData    => DMA0TXIRQ_GlitchData,
	OutSignalName => "DMA0TXIRQ",
	OutTemp       => DMA0TXIRQ_OUT,
	Paths         => (0 => (CPMDMA0LLCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => DMA1LLRSTENGINEACK,
	GlitchData    => DMA1LLRSTENGINEACK_GlitchData,
	OutSignalName => "DMA1LLRSTENGINEACK",
	OutTemp       => DMA1LLRSTENGINEACK_OUT,
	Paths         => (0 => (CPMDMA1LLCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => DMA1LLRXDSTRDYN,
	GlitchData    => DMA1LLRXDSTRDYN_GlitchData,
	OutSignalName => "DMA1LLRXDSTRDYN",
	OutTemp       => DMA1LLRXDSTRDYN_OUT,
	Paths         => (0 => (CPMDMA1LLCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => DMA1LLTXD(0),
	GlitchData    => DMA1LLTXD0_GlitchData,
	OutSignalName => "DMA1LLTXD(0)",
	OutTemp       => DMA1LLTXD_OUT(0),
	Paths         => (0 => (CPMDMA1LLCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => DMA1LLTXD(1),
	GlitchData    => DMA1LLTXD1_GlitchData,
	OutSignalName => "DMA1LLTXD(1)",
	OutTemp       => DMA1LLTXD_OUT(1),
	Paths         => (0 => (CPMDMA1LLCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => DMA1LLTXD(2),
	GlitchData    => DMA1LLTXD2_GlitchData,
	OutSignalName => "DMA1LLTXD(2)",
	OutTemp       => DMA1LLTXD_OUT(2),
	Paths         => (0 => (CPMDMA1LLCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => DMA1LLTXD(3),
	GlitchData    => DMA1LLTXD3_GlitchData,
	OutSignalName => "DMA1LLTXD(3)",
	OutTemp       => DMA1LLTXD_OUT(3),
	Paths         => (0 => (CPMDMA1LLCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => DMA1LLTXD(4),
	GlitchData    => DMA1LLTXD4_GlitchData,
	OutSignalName => "DMA1LLTXD(4)",
	OutTemp       => DMA1LLTXD_OUT(4),
	Paths         => (0 => (CPMDMA1LLCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => DMA1LLTXD(5),
	GlitchData    => DMA1LLTXD5_GlitchData,
	OutSignalName => "DMA1LLTXD(5)",
	OutTemp       => DMA1LLTXD_OUT(5),
	Paths         => (0 => (CPMDMA1LLCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => DMA1LLTXD(6),
	GlitchData    => DMA1LLTXD6_GlitchData,
	OutSignalName => "DMA1LLTXD(6)",
	OutTemp       => DMA1LLTXD_OUT(6),
	Paths         => (0 => (CPMDMA1LLCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => DMA1LLTXD(7),
	GlitchData    => DMA1LLTXD7_GlitchData,
	OutSignalName => "DMA1LLTXD(7)",
	OutTemp       => DMA1LLTXD_OUT(7),
	Paths         => (0 => (CPMDMA1LLCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => DMA1LLTXD(8),
	GlitchData    => DMA1LLTXD8_GlitchData,
	OutSignalName => "DMA1LLTXD(8)",
	OutTemp       => DMA1LLTXD_OUT(8),
	Paths         => (0 => (CPMDMA1LLCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => DMA1LLTXD(9),
	GlitchData    => DMA1LLTXD9_GlitchData,
	OutSignalName => "DMA1LLTXD(9)",
	OutTemp       => DMA1LLTXD_OUT(9),
	Paths         => (0 => (CPMDMA1LLCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => DMA1LLTXD(10),
	GlitchData    => DMA1LLTXD10_GlitchData,
	OutSignalName => "DMA1LLTXD(10)",
	OutTemp       => DMA1LLTXD_OUT(10),
	Paths         => (0 => (CPMDMA1LLCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => DMA1LLTXD(11),
	GlitchData    => DMA1LLTXD11_GlitchData,
	OutSignalName => "DMA1LLTXD(11)",
	OutTemp       => DMA1LLTXD_OUT(11),
	Paths         => (0 => (CPMDMA1LLCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => DMA1LLTXD(12),
	GlitchData    => DMA1LLTXD12_GlitchData,
	OutSignalName => "DMA1LLTXD(12)",
	OutTemp       => DMA1LLTXD_OUT(12),
	Paths         => (0 => (CPMDMA1LLCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => DMA1LLTXD(13),
	GlitchData    => DMA1LLTXD13_GlitchData,
	OutSignalName => "DMA1LLTXD(13)",
	OutTemp       => DMA1LLTXD_OUT(13),
	Paths         => (0 => (CPMDMA1LLCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => DMA1LLTXD(14),
	GlitchData    => DMA1LLTXD14_GlitchData,
	OutSignalName => "DMA1LLTXD(14)",
	OutTemp       => DMA1LLTXD_OUT(14),
	Paths         => (0 => (CPMDMA1LLCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => DMA1LLTXD(15),
	GlitchData    => DMA1LLTXD15_GlitchData,
	OutSignalName => "DMA1LLTXD(15)",
	OutTemp       => DMA1LLTXD_OUT(15),
	Paths         => (0 => (CPMDMA1LLCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => DMA1LLTXD(16),
	GlitchData    => DMA1LLTXD16_GlitchData,
	OutSignalName => "DMA1LLTXD(16)",
	OutTemp       => DMA1LLTXD_OUT(16),
	Paths         => (0 => (CPMDMA1LLCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => DMA1LLTXD(17),
	GlitchData    => DMA1LLTXD17_GlitchData,
	OutSignalName => "DMA1LLTXD(17)",
	OutTemp       => DMA1LLTXD_OUT(17),
	Paths         => (0 => (CPMDMA1LLCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => DMA1LLTXD(18),
	GlitchData    => DMA1LLTXD18_GlitchData,
	OutSignalName => "DMA1LLTXD(18)",
	OutTemp       => DMA1LLTXD_OUT(18),
	Paths         => (0 => (CPMDMA1LLCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => DMA1LLTXD(19),
	GlitchData    => DMA1LLTXD19_GlitchData,
	OutSignalName => "DMA1LLTXD(19)",
	OutTemp       => DMA1LLTXD_OUT(19),
	Paths         => (0 => (CPMDMA1LLCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => DMA1LLTXD(20),
	GlitchData    => DMA1LLTXD20_GlitchData,
	OutSignalName => "DMA1LLTXD(20)",
	OutTemp       => DMA1LLTXD_OUT(20),
	Paths         => (0 => (CPMDMA1LLCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => DMA1LLTXD(21),
	GlitchData    => DMA1LLTXD21_GlitchData,
	OutSignalName => "DMA1LLTXD(21)",
	OutTemp       => DMA1LLTXD_OUT(21),
	Paths         => (0 => (CPMDMA1LLCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => DMA1LLTXD(22),
	GlitchData    => DMA1LLTXD22_GlitchData,
	OutSignalName => "DMA1LLTXD(22)",
	OutTemp       => DMA1LLTXD_OUT(22),
	Paths         => (0 => (CPMDMA1LLCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => DMA1LLTXD(23),
	GlitchData    => DMA1LLTXD23_GlitchData,
	OutSignalName => "DMA1LLTXD(23)",
	OutTemp       => DMA1LLTXD_OUT(23),
	Paths         => (0 => (CPMDMA1LLCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => DMA1LLTXD(24),
	GlitchData    => DMA1LLTXD24_GlitchData,
	OutSignalName => "DMA1LLTXD(24)",
	OutTemp       => DMA1LLTXD_OUT(24),
	Paths         => (0 => (CPMDMA1LLCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => DMA1LLTXD(25),
	GlitchData    => DMA1LLTXD25_GlitchData,
	OutSignalName => "DMA1LLTXD(25)",
	OutTemp       => DMA1LLTXD_OUT(25),
	Paths         => (0 => (CPMDMA1LLCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => DMA1LLTXD(26),
	GlitchData    => DMA1LLTXD26_GlitchData,
	OutSignalName => "DMA1LLTXD(26)",
	OutTemp       => DMA1LLTXD_OUT(26),
	Paths         => (0 => (CPMDMA1LLCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => DMA1LLTXD(27),
	GlitchData    => DMA1LLTXD27_GlitchData,
	OutSignalName => "DMA1LLTXD(27)",
	OutTemp       => DMA1LLTXD_OUT(27),
	Paths         => (0 => (CPMDMA1LLCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => DMA1LLTXD(28),
	GlitchData    => DMA1LLTXD28_GlitchData,
	OutSignalName => "DMA1LLTXD(28)",
	OutTemp       => DMA1LLTXD_OUT(28),
	Paths         => (0 => (CPMDMA1LLCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => DMA1LLTXD(29),
	GlitchData    => DMA1LLTXD29_GlitchData,
	OutSignalName => "DMA1LLTXD(29)",
	OutTemp       => DMA1LLTXD_OUT(29),
	Paths         => (0 => (CPMDMA1LLCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => DMA1LLTXD(30),
	GlitchData    => DMA1LLTXD30_GlitchData,
	OutSignalName => "DMA1LLTXD(30)",
	OutTemp       => DMA1LLTXD_OUT(30),
	Paths         => (0 => (CPMDMA1LLCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => DMA1LLTXD(31),
	GlitchData    => DMA1LLTXD31_GlitchData,
	OutSignalName => "DMA1LLTXD(31)",
	OutTemp       => DMA1LLTXD_OUT(31),
	Paths         => (0 => (CPMDMA1LLCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => DMA1LLTXEOFN,
	GlitchData    => DMA1LLTXEOFN_GlitchData,
	OutSignalName => "DMA1LLTXEOFN",
	OutTemp       => DMA1LLTXEOFN_OUT,
	Paths         => (0 => (CPMDMA1LLCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => DMA1LLTXEOPN,
	GlitchData    => DMA1LLTXEOPN_GlitchData,
	OutSignalName => "DMA1LLTXEOPN",
	OutTemp       => DMA1LLTXEOPN_OUT,
	Paths         => (0 => (CPMDMA1LLCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => DMA1LLTXREM(0),
	GlitchData    => DMA1LLTXREM0_GlitchData,
	OutSignalName => "DMA1LLTXREM(0)",
	OutTemp       => DMA1LLTXREM_OUT(0),
	Paths         => (0 => (CPMDMA1LLCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => DMA1LLTXREM(1),
	GlitchData    => DMA1LLTXREM1_GlitchData,
	OutSignalName => "DMA1LLTXREM(1)",
	OutTemp       => DMA1LLTXREM_OUT(1),
	Paths         => (0 => (CPMDMA1LLCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => DMA1LLTXREM(2),
	GlitchData    => DMA1LLTXREM2_GlitchData,
	OutSignalName => "DMA1LLTXREM(2)",
	OutTemp       => DMA1LLTXREM_OUT(2),
	Paths         => (0 => (CPMDMA1LLCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => DMA1LLTXREM(3),
	GlitchData    => DMA1LLTXREM3_GlitchData,
	OutSignalName => "DMA1LLTXREM(3)",
	OutTemp       => DMA1LLTXREM_OUT(3),
	Paths         => (0 => (CPMDMA1LLCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => DMA1LLTXSOFN,
	GlitchData    => DMA1LLTXSOFN_GlitchData,
	OutSignalName => "DMA1LLTXSOFN",
	OutTemp       => DMA1LLTXSOFN_OUT,
	Paths         => (0 => (CPMDMA1LLCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => DMA1LLTXSOPN,
	GlitchData    => DMA1LLTXSOPN_GlitchData,
	OutSignalName => "DMA1LLTXSOPN",
	OutTemp       => DMA1LLTXSOPN_OUT,
	Paths         => (0 => (CPMDMA1LLCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => DMA1LLTXSRCRDYN,
	GlitchData    => DMA1LLTXSRCRDYN_GlitchData,
	OutSignalName => "DMA1LLTXSRCRDYN",
	OutTemp       => DMA1LLTXSRCRDYN_OUT,
	Paths         => (0 => (CPMDMA1LLCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => DMA1RXIRQ,
	GlitchData    => DMA1RXIRQ_GlitchData,
	OutSignalName => "DMA1RXIRQ",
	OutTemp       => DMA1RXIRQ_OUT,
	Paths         => (0 => (CPMDMA1LLCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => DMA1TXIRQ,
	GlitchData    => DMA1TXIRQ_GlitchData,
	OutSignalName => "DMA1TXIRQ",
	OutTemp       => DMA1TXIRQ_OUT,
	Paths         => (0 => (CPMDMA1LLCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => DMA2LLRSTENGINEACK,
	GlitchData    => DMA2LLRSTENGINEACK_GlitchData,
	OutSignalName => "DMA2LLRSTENGINEACK",
	OutTemp       => DMA2LLRSTENGINEACK_OUT,
	Paths         => (0 => (CPMDMA2LLCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => DMA2LLRXDSTRDYN,
	GlitchData    => DMA2LLRXDSTRDYN_GlitchData,
	OutSignalName => "DMA2LLRXDSTRDYN",
	OutTemp       => DMA2LLRXDSTRDYN_OUT,
	Paths         => (0 => (CPMDMA2LLCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => DMA2LLTXD(0),
	GlitchData    => DMA2LLTXD0_GlitchData,
	OutSignalName => "DMA2LLTXD(0)",
	OutTemp       => DMA2LLTXD_OUT(0),
	Paths         => (0 => (CPMDMA2LLCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => DMA2LLTXD(1),
	GlitchData    => DMA2LLTXD1_GlitchData,
	OutSignalName => "DMA2LLTXD(1)",
	OutTemp       => DMA2LLTXD_OUT(1),
	Paths         => (0 => (CPMDMA2LLCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => DMA2LLTXD(2),
	GlitchData    => DMA2LLTXD2_GlitchData,
	OutSignalName => "DMA2LLTXD(2)",
	OutTemp       => DMA2LLTXD_OUT(2),
	Paths         => (0 => (CPMDMA2LLCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => DMA2LLTXD(3),
	GlitchData    => DMA2LLTXD3_GlitchData,
	OutSignalName => "DMA2LLTXD(3)",
	OutTemp       => DMA2LLTXD_OUT(3),
	Paths         => (0 => (CPMDMA2LLCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => DMA2LLTXD(4),
	GlitchData    => DMA2LLTXD4_GlitchData,
	OutSignalName => "DMA2LLTXD(4)",
	OutTemp       => DMA2LLTXD_OUT(4),
	Paths         => (0 => (CPMDMA2LLCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => DMA2LLTXD(5),
	GlitchData    => DMA2LLTXD5_GlitchData,
	OutSignalName => "DMA2LLTXD(5)",
	OutTemp       => DMA2LLTXD_OUT(5),
	Paths         => (0 => (CPMDMA2LLCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => DMA2LLTXD(6),
	GlitchData    => DMA2LLTXD6_GlitchData,
	OutSignalName => "DMA2LLTXD(6)",
	OutTemp       => DMA2LLTXD_OUT(6),
	Paths         => (0 => (CPMDMA2LLCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => DMA2LLTXD(7),
	GlitchData    => DMA2LLTXD7_GlitchData,
	OutSignalName => "DMA2LLTXD(7)",
	OutTemp       => DMA2LLTXD_OUT(7),
	Paths         => (0 => (CPMDMA2LLCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => DMA2LLTXD(8),
	GlitchData    => DMA2LLTXD8_GlitchData,
	OutSignalName => "DMA2LLTXD(8)",
	OutTemp       => DMA2LLTXD_OUT(8),
	Paths         => (0 => (CPMDMA2LLCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => DMA2LLTXD(9),
	GlitchData    => DMA2LLTXD9_GlitchData,
	OutSignalName => "DMA2LLTXD(9)",
	OutTemp       => DMA2LLTXD_OUT(9),
	Paths         => (0 => (CPMDMA2LLCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => DMA2LLTXD(10),
	GlitchData    => DMA2LLTXD10_GlitchData,
	OutSignalName => "DMA2LLTXD(10)",
	OutTemp       => DMA2LLTXD_OUT(10),
	Paths         => (0 => (CPMDMA2LLCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => DMA2LLTXD(11),
	GlitchData    => DMA2LLTXD11_GlitchData,
	OutSignalName => "DMA2LLTXD(11)",
	OutTemp       => DMA2LLTXD_OUT(11),
	Paths         => (0 => (CPMDMA2LLCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => DMA2LLTXD(12),
	GlitchData    => DMA2LLTXD12_GlitchData,
	OutSignalName => "DMA2LLTXD(12)",
	OutTemp       => DMA2LLTXD_OUT(12),
	Paths         => (0 => (CPMDMA2LLCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => DMA2LLTXD(13),
	GlitchData    => DMA2LLTXD13_GlitchData,
	OutSignalName => "DMA2LLTXD(13)",
	OutTemp       => DMA2LLTXD_OUT(13),
	Paths         => (0 => (CPMDMA2LLCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => DMA2LLTXD(14),
	GlitchData    => DMA2LLTXD14_GlitchData,
	OutSignalName => "DMA2LLTXD(14)",
	OutTemp       => DMA2LLTXD_OUT(14),
	Paths         => (0 => (CPMDMA2LLCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => DMA2LLTXD(15),
	GlitchData    => DMA2LLTXD15_GlitchData,
	OutSignalName => "DMA2LLTXD(15)",
	OutTemp       => DMA2LLTXD_OUT(15),
	Paths         => (0 => (CPMDMA2LLCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => DMA2LLTXD(16),
	GlitchData    => DMA2LLTXD16_GlitchData,
	OutSignalName => "DMA2LLTXD(16)",
	OutTemp       => DMA2LLTXD_OUT(16),
	Paths         => (0 => (CPMDMA2LLCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => DMA2LLTXD(17),
	GlitchData    => DMA2LLTXD17_GlitchData,
	OutSignalName => "DMA2LLTXD(17)",
	OutTemp       => DMA2LLTXD_OUT(17),
	Paths         => (0 => (CPMDMA2LLCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => DMA2LLTXD(18),
	GlitchData    => DMA2LLTXD18_GlitchData,
	OutSignalName => "DMA2LLTXD(18)",
	OutTemp       => DMA2LLTXD_OUT(18),
	Paths         => (0 => (CPMDMA2LLCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => DMA2LLTXD(19),
	GlitchData    => DMA2LLTXD19_GlitchData,
	OutSignalName => "DMA2LLTXD(19)",
	OutTemp       => DMA2LLTXD_OUT(19),
	Paths         => (0 => (CPMDMA2LLCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => DMA2LLTXD(20),
	GlitchData    => DMA2LLTXD20_GlitchData,
	OutSignalName => "DMA2LLTXD(20)",
	OutTemp       => DMA2LLTXD_OUT(20),
	Paths         => (0 => (CPMDMA2LLCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => DMA2LLTXD(21),
	GlitchData    => DMA2LLTXD21_GlitchData,
	OutSignalName => "DMA2LLTXD(21)",
	OutTemp       => DMA2LLTXD_OUT(21),
	Paths         => (0 => (CPMDMA2LLCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => DMA2LLTXD(22),
	GlitchData    => DMA2LLTXD22_GlitchData,
	OutSignalName => "DMA2LLTXD(22)",
	OutTemp       => DMA2LLTXD_OUT(22),
	Paths         => (0 => (CPMDMA2LLCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => DMA2LLTXD(23),
	GlitchData    => DMA2LLTXD23_GlitchData,
	OutSignalName => "DMA2LLTXD(23)",
	OutTemp       => DMA2LLTXD_OUT(23),
	Paths         => (0 => (CPMDMA2LLCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => DMA2LLTXD(24),
	GlitchData    => DMA2LLTXD24_GlitchData,
	OutSignalName => "DMA2LLTXD(24)",
	OutTemp       => DMA2LLTXD_OUT(24),
	Paths         => (0 => (CPMDMA2LLCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => DMA2LLTXD(25),
	GlitchData    => DMA2LLTXD25_GlitchData,
	OutSignalName => "DMA2LLTXD(25)",
	OutTemp       => DMA2LLTXD_OUT(25),
	Paths         => (0 => (CPMDMA2LLCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => DMA2LLTXD(26),
	GlitchData    => DMA2LLTXD26_GlitchData,
	OutSignalName => "DMA2LLTXD(26)",
	OutTemp       => DMA2LLTXD_OUT(26),
	Paths         => (0 => (CPMDMA2LLCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => DMA2LLTXD(27),
	GlitchData    => DMA2LLTXD27_GlitchData,
	OutSignalName => "DMA2LLTXD(27)",
	OutTemp       => DMA2LLTXD_OUT(27),
	Paths         => (0 => (CPMDMA2LLCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => DMA2LLTXD(28),
	GlitchData    => DMA2LLTXD28_GlitchData,
	OutSignalName => "DMA2LLTXD(28)",
	OutTemp       => DMA2LLTXD_OUT(28),
	Paths         => (0 => (CPMDMA2LLCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => DMA2LLTXD(29),
	GlitchData    => DMA2LLTXD29_GlitchData,
	OutSignalName => "DMA2LLTXD(29)",
	OutTemp       => DMA2LLTXD_OUT(29),
	Paths         => (0 => (CPMDMA2LLCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => DMA2LLTXD(30),
	GlitchData    => DMA2LLTXD30_GlitchData,
	OutSignalName => "DMA2LLTXD(30)",
	OutTemp       => DMA2LLTXD_OUT(30),
	Paths         => (0 => (CPMDMA2LLCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => DMA2LLTXD(31),
	GlitchData    => DMA2LLTXD31_GlitchData,
	OutSignalName => "DMA2LLTXD(31)",
	OutTemp       => DMA2LLTXD_OUT(31),
	Paths         => (0 => (CPMDMA2LLCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => DMA2LLTXEOFN,
	GlitchData    => DMA2LLTXEOFN_GlitchData,
	OutSignalName => "DMA2LLTXEOFN",
	OutTemp       => DMA2LLTXEOFN_OUT,
	Paths         => (0 => (CPMDMA2LLCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => DMA2LLTXEOPN,
	GlitchData    => DMA2LLTXEOPN_GlitchData,
	OutSignalName => "DMA2LLTXEOPN",
	OutTemp       => DMA2LLTXEOPN_OUT,
	Paths         => (0 => (CPMDMA2LLCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => DMA2LLTXREM(0),
	GlitchData    => DMA2LLTXREM0_GlitchData,
	OutSignalName => "DMA2LLTXREM(0)",
	OutTemp       => DMA2LLTXREM_OUT(0),
	Paths         => (0 => (CPMDMA2LLCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => DMA2LLTXREM(1),
	GlitchData    => DMA2LLTXREM1_GlitchData,
	OutSignalName => "DMA2LLTXREM(1)",
	OutTemp       => DMA2LLTXREM_OUT(1),
	Paths         => (0 => (CPMDMA2LLCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => DMA2LLTXREM(2),
	GlitchData    => DMA2LLTXREM2_GlitchData,
	OutSignalName => "DMA2LLTXREM(2)",
	OutTemp       => DMA2LLTXREM_OUT(2),
	Paths         => (0 => (CPMDMA2LLCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => DMA2LLTXREM(3),
	GlitchData    => DMA2LLTXREM3_GlitchData,
	OutSignalName => "DMA2LLTXREM(3)",
	OutTemp       => DMA2LLTXREM_OUT(3),
	Paths         => (0 => (CPMDMA2LLCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => DMA2LLTXSOFN,
	GlitchData    => DMA2LLTXSOFN_GlitchData,
	OutSignalName => "DMA2LLTXSOFN",
	OutTemp       => DMA2LLTXSOFN_OUT,
	Paths         => (0 => (CPMDMA2LLCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => DMA2LLTXSOPN,
	GlitchData    => DMA2LLTXSOPN_GlitchData,
	OutSignalName => "DMA2LLTXSOPN",
	OutTemp       => DMA2LLTXSOPN_OUT,
	Paths         => (0 => (CPMDMA2LLCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => DMA2LLTXSRCRDYN,
	GlitchData    => DMA2LLTXSRCRDYN_GlitchData,
	OutSignalName => "DMA2LLTXSRCRDYN",
	OutTemp       => DMA2LLTXSRCRDYN_OUT,
	Paths         => (0 => (CPMDMA2LLCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => DMA2RXIRQ,
	GlitchData    => DMA2RXIRQ_GlitchData,
	OutSignalName => "DMA2RXIRQ",
	OutTemp       => DMA2RXIRQ_OUT,
	Paths         => (0 => (CPMDMA2LLCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => DMA2TXIRQ,
	GlitchData    => DMA2TXIRQ_GlitchData,
	OutSignalName => "DMA2TXIRQ",
	OutTemp       => DMA2TXIRQ_OUT,
	Paths         => (0 => (CPMDMA2LLCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => DMA3LLRSTENGINEACK,
	GlitchData    => DMA3LLRSTENGINEACK_GlitchData,
	OutSignalName => "DMA3LLRSTENGINEACK",
	OutTemp       => DMA3LLRSTENGINEACK_OUT,
	Paths         => (0 => (CPMDMA3LLCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => DMA3LLRXDSTRDYN,
	GlitchData    => DMA3LLRXDSTRDYN_GlitchData,
	OutSignalName => "DMA3LLRXDSTRDYN",
	OutTemp       => DMA3LLRXDSTRDYN_OUT,
	Paths         => (0 => (CPMDMA3LLCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => DMA3LLTXD(0),
	GlitchData    => DMA3LLTXD0_GlitchData,
	OutSignalName => "DMA3LLTXD(0)",
	OutTemp       => DMA3LLTXD_OUT(0),
	Paths         => (0 => (CPMDMA3LLCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => DMA3LLTXD(1),
	GlitchData    => DMA3LLTXD1_GlitchData,
	OutSignalName => "DMA3LLTXD(1)",
	OutTemp       => DMA3LLTXD_OUT(1),
	Paths         => (0 => (CPMDMA3LLCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => DMA3LLTXD(2),
	GlitchData    => DMA3LLTXD2_GlitchData,
	OutSignalName => "DMA3LLTXD(2)",
	OutTemp       => DMA3LLTXD_OUT(2),
	Paths         => (0 => (CPMDMA3LLCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => DMA3LLTXD(3),
	GlitchData    => DMA3LLTXD3_GlitchData,
	OutSignalName => "DMA3LLTXD(3)",
	OutTemp       => DMA3LLTXD_OUT(3),
	Paths         => (0 => (CPMDMA3LLCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => DMA3LLTXD(4),
	GlitchData    => DMA3LLTXD4_GlitchData,
	OutSignalName => "DMA3LLTXD(4)",
	OutTemp       => DMA3LLTXD_OUT(4),
	Paths         => (0 => (CPMDMA3LLCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => DMA3LLTXD(5),
	GlitchData    => DMA3LLTXD5_GlitchData,
	OutSignalName => "DMA3LLTXD(5)",
	OutTemp       => DMA3LLTXD_OUT(5),
	Paths         => (0 => (CPMDMA3LLCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => DMA3LLTXD(6),
	GlitchData    => DMA3LLTXD6_GlitchData,
	OutSignalName => "DMA3LLTXD(6)",
	OutTemp       => DMA3LLTXD_OUT(6),
	Paths         => (0 => (CPMDMA3LLCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => DMA3LLTXD(7),
	GlitchData    => DMA3LLTXD7_GlitchData,
	OutSignalName => "DMA3LLTXD(7)",
	OutTemp       => DMA3LLTXD_OUT(7),
	Paths         => (0 => (CPMDMA3LLCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => DMA3LLTXD(8),
	GlitchData    => DMA3LLTXD8_GlitchData,
	OutSignalName => "DMA3LLTXD(8)",
	OutTemp       => DMA3LLTXD_OUT(8),
	Paths         => (0 => (CPMDMA3LLCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => DMA3LLTXD(9),
	GlitchData    => DMA3LLTXD9_GlitchData,
	OutSignalName => "DMA3LLTXD(9)",
	OutTemp       => DMA3LLTXD_OUT(9),
	Paths         => (0 => (CPMDMA3LLCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => DMA3LLTXD(10),
	GlitchData    => DMA3LLTXD10_GlitchData,
	OutSignalName => "DMA3LLTXD(10)",
	OutTemp       => DMA3LLTXD_OUT(10),
	Paths         => (0 => (CPMDMA3LLCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => DMA3LLTXD(11),
	GlitchData    => DMA3LLTXD11_GlitchData,
	OutSignalName => "DMA3LLTXD(11)",
	OutTemp       => DMA3LLTXD_OUT(11),
	Paths         => (0 => (CPMDMA3LLCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => DMA3LLTXD(12),
	GlitchData    => DMA3LLTXD12_GlitchData,
	OutSignalName => "DMA3LLTXD(12)",
	OutTemp       => DMA3LLTXD_OUT(12),
	Paths         => (0 => (CPMDMA3LLCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => DMA3LLTXD(13),
	GlitchData    => DMA3LLTXD13_GlitchData,
	OutSignalName => "DMA3LLTXD(13)",
	OutTemp       => DMA3LLTXD_OUT(13),
	Paths         => (0 => (CPMDMA3LLCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => DMA3LLTXD(14),
	GlitchData    => DMA3LLTXD14_GlitchData,
	OutSignalName => "DMA3LLTXD(14)",
	OutTemp       => DMA3LLTXD_OUT(14),
	Paths         => (0 => (CPMDMA3LLCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => DMA3LLTXD(15),
	GlitchData    => DMA3LLTXD15_GlitchData,
	OutSignalName => "DMA3LLTXD(15)",
	OutTemp       => DMA3LLTXD_OUT(15),
	Paths         => (0 => (CPMDMA3LLCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => DMA3LLTXD(16),
	GlitchData    => DMA3LLTXD16_GlitchData,
	OutSignalName => "DMA3LLTXD(16)",
	OutTemp       => DMA3LLTXD_OUT(16),
	Paths         => (0 => (CPMDMA3LLCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => DMA3LLTXD(17),
	GlitchData    => DMA3LLTXD17_GlitchData,
	OutSignalName => "DMA3LLTXD(17)",
	OutTemp       => DMA3LLTXD_OUT(17),
	Paths         => (0 => (CPMDMA3LLCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => DMA3LLTXD(18),
	GlitchData    => DMA3LLTXD18_GlitchData,
	OutSignalName => "DMA3LLTXD(18)",
	OutTemp       => DMA3LLTXD_OUT(18),
	Paths         => (0 => (CPMDMA3LLCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => DMA3LLTXD(19),
	GlitchData    => DMA3LLTXD19_GlitchData,
	OutSignalName => "DMA3LLTXD(19)",
	OutTemp       => DMA3LLTXD_OUT(19),
	Paths         => (0 => (CPMDMA3LLCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => DMA3LLTXD(20),
	GlitchData    => DMA3LLTXD20_GlitchData,
	OutSignalName => "DMA3LLTXD(20)",
	OutTemp       => DMA3LLTXD_OUT(20),
	Paths         => (0 => (CPMDMA3LLCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => DMA3LLTXD(21),
	GlitchData    => DMA3LLTXD21_GlitchData,
	OutSignalName => "DMA3LLTXD(21)",
	OutTemp       => DMA3LLTXD_OUT(21),
	Paths         => (0 => (CPMDMA3LLCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => DMA3LLTXD(22),
	GlitchData    => DMA3LLTXD22_GlitchData,
	OutSignalName => "DMA3LLTXD(22)",
	OutTemp       => DMA3LLTXD_OUT(22),
	Paths         => (0 => (CPMDMA3LLCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => DMA3LLTXD(23),
	GlitchData    => DMA3LLTXD23_GlitchData,
	OutSignalName => "DMA3LLTXD(23)",
	OutTemp       => DMA3LLTXD_OUT(23),
	Paths         => (0 => (CPMDMA3LLCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => DMA3LLTXD(24),
	GlitchData    => DMA3LLTXD24_GlitchData,
	OutSignalName => "DMA3LLTXD(24)",
	OutTemp       => DMA3LLTXD_OUT(24),
	Paths         => (0 => (CPMDMA3LLCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => DMA3LLTXD(25),
	GlitchData    => DMA3LLTXD25_GlitchData,
	OutSignalName => "DMA3LLTXD(25)",
	OutTemp       => DMA3LLTXD_OUT(25),
	Paths         => (0 => (CPMDMA3LLCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => DMA3LLTXD(26),
	GlitchData    => DMA3LLTXD26_GlitchData,
	OutSignalName => "DMA3LLTXD(26)",
	OutTemp       => DMA3LLTXD_OUT(26),
	Paths         => (0 => (CPMDMA3LLCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => DMA3LLTXD(27),
	GlitchData    => DMA3LLTXD27_GlitchData,
	OutSignalName => "DMA3LLTXD(27)",
	OutTemp       => DMA3LLTXD_OUT(27),
	Paths         => (0 => (CPMDMA3LLCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => DMA3LLTXD(28),
	GlitchData    => DMA3LLTXD28_GlitchData,
	OutSignalName => "DMA3LLTXD(28)",
	OutTemp       => DMA3LLTXD_OUT(28),
	Paths         => (0 => (CPMDMA3LLCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => DMA3LLTXD(29),
	GlitchData    => DMA3LLTXD29_GlitchData,
	OutSignalName => "DMA3LLTXD(29)",
	OutTemp       => DMA3LLTXD_OUT(29),
	Paths         => (0 => (CPMDMA3LLCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => DMA3LLTXD(30),
	GlitchData    => DMA3LLTXD30_GlitchData,
	OutSignalName => "DMA3LLTXD(30)",
	OutTemp       => DMA3LLTXD_OUT(30),
	Paths         => (0 => (CPMDMA3LLCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => DMA3LLTXD(31),
	GlitchData    => DMA3LLTXD31_GlitchData,
	OutSignalName => "DMA3LLTXD(31)",
	OutTemp       => DMA3LLTXD_OUT(31),
	Paths         => (0 => (CPMDMA3LLCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => DMA3LLTXEOFN,
	GlitchData    => DMA3LLTXEOFN_GlitchData,
	OutSignalName => "DMA3LLTXEOFN",
	OutTemp       => DMA3LLTXEOFN_OUT,
	Paths         => (0 => (CPMDMA3LLCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => DMA3LLTXEOPN,
	GlitchData    => DMA3LLTXEOPN_GlitchData,
	OutSignalName => "DMA3LLTXEOPN",
	OutTemp       => DMA3LLTXEOPN_OUT,
	Paths         => (0 => (CPMDMA3LLCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => DMA3LLTXREM(0),
	GlitchData    => DMA3LLTXREM0_GlitchData,
	OutSignalName => "DMA3LLTXREM(0)",
	OutTemp       => DMA3LLTXREM_OUT(0),
	Paths         => (0 => (CPMDMA3LLCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => DMA3LLTXREM(1),
	GlitchData    => DMA3LLTXREM1_GlitchData,
	OutSignalName => "DMA3LLTXREM(1)",
	OutTemp       => DMA3LLTXREM_OUT(1),
	Paths         => (0 => (CPMDMA3LLCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => DMA3LLTXREM(2),
	GlitchData    => DMA3LLTXREM2_GlitchData,
	OutSignalName => "DMA3LLTXREM(2)",
	OutTemp       => DMA3LLTXREM_OUT(2),
	Paths         => (0 => (CPMDMA3LLCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => DMA3LLTXREM(3),
	GlitchData    => DMA3LLTXREM3_GlitchData,
	OutSignalName => "DMA3LLTXREM(3)",
	OutTemp       => DMA3LLTXREM_OUT(3),
	Paths         => (0 => (CPMDMA3LLCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => DMA3LLTXSOFN,
	GlitchData    => DMA3LLTXSOFN_GlitchData,
	OutSignalName => "DMA3LLTXSOFN",
	OutTemp       => DMA3LLTXSOFN_OUT,
	Paths         => (0 => (CPMDMA3LLCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => DMA3LLTXSOPN,
	GlitchData    => DMA3LLTXSOPN_GlitchData,
	OutSignalName => "DMA3LLTXSOPN",
	OutTemp       => DMA3LLTXSOPN_OUT,
	Paths         => (0 => (CPMDMA3LLCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => DMA3LLTXSRCRDYN,
	GlitchData    => DMA3LLTXSRCRDYN_GlitchData,
	OutSignalName => "DMA3LLTXSRCRDYN",
	OutTemp       => DMA3LLTXSRCRDYN_OUT,
	Paths         => (0 => (CPMDMA3LLCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => DMA3RXIRQ,
	GlitchData    => DMA3RXIRQ_GlitchData,
	OutSignalName => "DMA3RXIRQ",
	OutTemp       => DMA3RXIRQ_OUT,
	Paths         => (0 => (CPMDMA3LLCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => DMA3TXIRQ,
	GlitchData    => DMA3TXIRQ_GlitchData,
	OutSignalName => "DMA3TXIRQ",
	OutTemp       => DMA3TXIRQ_OUT,
	Paths         => (0 => (CPMDMA3LLCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCDMDCRABUS(0),
	GlitchData    => PPCDMDCRABUS0_GlitchData,
	OutSignalName => "PPCDMDCRABUS(0)",
	OutTemp       => PPCDMDCRABUS_OUT(0),
	Paths         => (0 => (CPMDCRCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCDMDCRABUS(1),
	GlitchData    => PPCDMDCRABUS1_GlitchData,
	OutSignalName => "PPCDMDCRABUS(1)",
	OutTemp       => PPCDMDCRABUS_OUT(1),
	Paths         => (0 => (CPMDCRCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCDMDCRABUS(2),
	GlitchData    => PPCDMDCRABUS2_GlitchData,
	OutSignalName => "PPCDMDCRABUS(2)",
	OutTemp       => PPCDMDCRABUS_OUT(2),
	Paths         => (0 => (CPMDCRCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCDMDCRABUS(3),
	GlitchData    => PPCDMDCRABUS3_GlitchData,
	OutSignalName => "PPCDMDCRABUS(3)",
	OutTemp       => PPCDMDCRABUS_OUT(3),
	Paths         => (0 => (CPMDCRCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCDMDCRABUS(4),
	GlitchData    => PPCDMDCRABUS4_GlitchData,
	OutSignalName => "PPCDMDCRABUS(4)",
	OutTemp       => PPCDMDCRABUS_OUT(4),
	Paths         => (0 => (CPMDCRCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCDMDCRABUS(5),
	GlitchData    => PPCDMDCRABUS5_GlitchData,
	OutSignalName => "PPCDMDCRABUS(5)",
	OutTemp       => PPCDMDCRABUS_OUT(5),
	Paths         => (0 => (CPMDCRCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCDMDCRABUS(6),
	GlitchData    => PPCDMDCRABUS6_GlitchData,
	OutSignalName => "PPCDMDCRABUS(6)",
	OutTemp       => PPCDMDCRABUS_OUT(6),
	Paths         => (0 => (CPMDCRCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCDMDCRABUS(7),
	GlitchData    => PPCDMDCRABUS7_GlitchData,
	OutSignalName => "PPCDMDCRABUS(7)",
	OutTemp       => PPCDMDCRABUS_OUT(7),
	Paths         => (0 => (CPMDCRCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCDMDCRABUS(8),
	GlitchData    => PPCDMDCRABUS8_GlitchData,
	OutSignalName => "PPCDMDCRABUS(8)",
	OutTemp       => PPCDMDCRABUS_OUT(8),
	Paths         => (0 => (CPMDCRCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCDMDCRABUS(9),
	GlitchData    => PPCDMDCRABUS9_GlitchData,
	OutSignalName => "PPCDMDCRABUS(9)",
	OutTemp       => PPCDMDCRABUS_OUT(9),
	Paths         => (0 => (CPMDCRCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCDMDCRDBUSOUT(0),
	GlitchData    => PPCDMDCRDBUSOUT0_GlitchData,
	OutSignalName => "PPCDMDCRDBUSOUT(0)",
	OutTemp       => PPCDMDCRDBUSOUT_OUT(0),
	Paths         => (0 => (CPMDCRCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCDMDCRDBUSOUT(1),
	GlitchData    => PPCDMDCRDBUSOUT1_GlitchData,
	OutSignalName => "PPCDMDCRDBUSOUT(1)",
	OutTemp       => PPCDMDCRDBUSOUT_OUT(1),
	Paths         => (0 => (CPMDCRCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCDMDCRDBUSOUT(2),
	GlitchData    => PPCDMDCRDBUSOUT2_GlitchData,
	OutSignalName => "PPCDMDCRDBUSOUT(2)",
	OutTemp       => PPCDMDCRDBUSOUT_OUT(2),
	Paths         => (0 => (CPMDCRCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCDMDCRDBUSOUT(3),
	GlitchData    => PPCDMDCRDBUSOUT3_GlitchData,
	OutSignalName => "PPCDMDCRDBUSOUT(3)",
	OutTemp       => PPCDMDCRDBUSOUT_OUT(3),
	Paths         => (0 => (CPMDCRCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCDMDCRDBUSOUT(4),
	GlitchData    => PPCDMDCRDBUSOUT4_GlitchData,
	OutSignalName => "PPCDMDCRDBUSOUT(4)",
	OutTemp       => PPCDMDCRDBUSOUT_OUT(4),
	Paths         => (0 => (CPMDCRCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCDMDCRDBUSOUT(5),
	GlitchData    => PPCDMDCRDBUSOUT5_GlitchData,
	OutSignalName => "PPCDMDCRDBUSOUT(5)",
	OutTemp       => PPCDMDCRDBUSOUT_OUT(5),
	Paths         => (0 => (CPMDCRCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCDMDCRDBUSOUT(6),
	GlitchData    => PPCDMDCRDBUSOUT6_GlitchData,
	OutSignalName => "PPCDMDCRDBUSOUT(6)",
	OutTemp       => PPCDMDCRDBUSOUT_OUT(6),
	Paths         => (0 => (CPMDCRCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCDMDCRDBUSOUT(7),
	GlitchData    => PPCDMDCRDBUSOUT7_GlitchData,
	OutSignalName => "PPCDMDCRDBUSOUT(7)",
	OutTemp       => PPCDMDCRDBUSOUT_OUT(7),
	Paths         => (0 => (CPMDCRCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCDMDCRDBUSOUT(8),
	GlitchData    => PPCDMDCRDBUSOUT8_GlitchData,
	OutSignalName => "PPCDMDCRDBUSOUT(8)",
	OutTemp       => PPCDMDCRDBUSOUT_OUT(8),
	Paths         => (0 => (CPMDCRCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCDMDCRDBUSOUT(9),
	GlitchData    => PPCDMDCRDBUSOUT9_GlitchData,
	OutSignalName => "PPCDMDCRDBUSOUT(9)",
	OutTemp       => PPCDMDCRDBUSOUT_OUT(9),
	Paths         => (0 => (CPMDCRCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCDMDCRDBUSOUT(10),
	GlitchData    => PPCDMDCRDBUSOUT10_GlitchData,
	OutSignalName => "PPCDMDCRDBUSOUT(10)",
	OutTemp       => PPCDMDCRDBUSOUT_OUT(10),
	Paths         => (0 => (CPMDCRCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCDMDCRDBUSOUT(11),
	GlitchData    => PPCDMDCRDBUSOUT11_GlitchData,
	OutSignalName => "PPCDMDCRDBUSOUT(11)",
	OutTemp       => PPCDMDCRDBUSOUT_OUT(11),
	Paths         => (0 => (CPMDCRCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCDMDCRDBUSOUT(12),
	GlitchData    => PPCDMDCRDBUSOUT12_GlitchData,
	OutSignalName => "PPCDMDCRDBUSOUT(12)",
	OutTemp       => PPCDMDCRDBUSOUT_OUT(12),
	Paths         => (0 => (CPMDCRCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCDMDCRDBUSOUT(13),
	GlitchData    => PPCDMDCRDBUSOUT13_GlitchData,
	OutSignalName => "PPCDMDCRDBUSOUT(13)",
	OutTemp       => PPCDMDCRDBUSOUT_OUT(13),
	Paths         => (0 => (CPMDCRCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCDMDCRDBUSOUT(14),
	GlitchData    => PPCDMDCRDBUSOUT14_GlitchData,
	OutSignalName => "PPCDMDCRDBUSOUT(14)",
	OutTemp       => PPCDMDCRDBUSOUT_OUT(14),
	Paths         => (0 => (CPMDCRCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCDMDCRDBUSOUT(15),
	GlitchData    => PPCDMDCRDBUSOUT15_GlitchData,
	OutSignalName => "PPCDMDCRDBUSOUT(15)",
	OutTemp       => PPCDMDCRDBUSOUT_OUT(15),
	Paths         => (0 => (CPMDCRCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCDMDCRDBUSOUT(16),
	GlitchData    => PPCDMDCRDBUSOUT16_GlitchData,
	OutSignalName => "PPCDMDCRDBUSOUT(16)",
	OutTemp       => PPCDMDCRDBUSOUT_OUT(16),
	Paths         => (0 => (CPMDCRCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCDMDCRDBUSOUT(17),
	GlitchData    => PPCDMDCRDBUSOUT17_GlitchData,
	OutSignalName => "PPCDMDCRDBUSOUT(17)",
	OutTemp       => PPCDMDCRDBUSOUT_OUT(17),
	Paths         => (0 => (CPMDCRCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCDMDCRDBUSOUT(18),
	GlitchData    => PPCDMDCRDBUSOUT18_GlitchData,
	OutSignalName => "PPCDMDCRDBUSOUT(18)",
	OutTemp       => PPCDMDCRDBUSOUT_OUT(18),
	Paths         => (0 => (CPMDCRCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCDMDCRDBUSOUT(19),
	GlitchData    => PPCDMDCRDBUSOUT19_GlitchData,
	OutSignalName => "PPCDMDCRDBUSOUT(19)",
	OutTemp       => PPCDMDCRDBUSOUT_OUT(19),
	Paths         => (0 => (CPMDCRCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCDMDCRDBUSOUT(20),
	GlitchData    => PPCDMDCRDBUSOUT20_GlitchData,
	OutSignalName => "PPCDMDCRDBUSOUT(20)",
	OutTemp       => PPCDMDCRDBUSOUT_OUT(20),
	Paths         => (0 => (CPMDCRCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCDMDCRDBUSOUT(21),
	GlitchData    => PPCDMDCRDBUSOUT21_GlitchData,
	OutSignalName => "PPCDMDCRDBUSOUT(21)",
	OutTemp       => PPCDMDCRDBUSOUT_OUT(21),
	Paths         => (0 => (CPMDCRCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCDMDCRDBUSOUT(22),
	GlitchData    => PPCDMDCRDBUSOUT22_GlitchData,
	OutSignalName => "PPCDMDCRDBUSOUT(22)",
	OutTemp       => PPCDMDCRDBUSOUT_OUT(22),
	Paths         => (0 => (CPMDCRCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCDMDCRDBUSOUT(23),
	GlitchData    => PPCDMDCRDBUSOUT23_GlitchData,
	OutSignalName => "PPCDMDCRDBUSOUT(23)",
	OutTemp       => PPCDMDCRDBUSOUT_OUT(23),
	Paths         => (0 => (CPMDCRCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCDMDCRDBUSOUT(24),
	GlitchData    => PPCDMDCRDBUSOUT24_GlitchData,
	OutSignalName => "PPCDMDCRDBUSOUT(24)",
	OutTemp       => PPCDMDCRDBUSOUT_OUT(24),
	Paths         => (0 => (CPMDCRCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCDMDCRDBUSOUT(25),
	GlitchData    => PPCDMDCRDBUSOUT25_GlitchData,
	OutSignalName => "PPCDMDCRDBUSOUT(25)",
	OutTemp       => PPCDMDCRDBUSOUT_OUT(25),
	Paths         => (0 => (CPMDCRCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCDMDCRDBUSOUT(26),
	GlitchData    => PPCDMDCRDBUSOUT26_GlitchData,
	OutSignalName => "PPCDMDCRDBUSOUT(26)",
	OutTemp       => PPCDMDCRDBUSOUT_OUT(26),
	Paths         => (0 => (CPMDCRCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCDMDCRDBUSOUT(27),
	GlitchData    => PPCDMDCRDBUSOUT27_GlitchData,
	OutSignalName => "PPCDMDCRDBUSOUT(27)",
	OutTemp       => PPCDMDCRDBUSOUT_OUT(27),
	Paths         => (0 => (CPMDCRCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCDMDCRDBUSOUT(28),
	GlitchData    => PPCDMDCRDBUSOUT28_GlitchData,
	OutSignalName => "PPCDMDCRDBUSOUT(28)",
	OutTemp       => PPCDMDCRDBUSOUT_OUT(28),
	Paths         => (0 => (CPMDCRCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCDMDCRDBUSOUT(29),
	GlitchData    => PPCDMDCRDBUSOUT29_GlitchData,
	OutSignalName => "PPCDMDCRDBUSOUT(29)",
	OutTemp       => PPCDMDCRDBUSOUT_OUT(29),
	Paths         => (0 => (CPMDCRCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCDMDCRDBUSOUT(30),
	GlitchData    => PPCDMDCRDBUSOUT30_GlitchData,
	OutSignalName => "PPCDMDCRDBUSOUT(30)",
	OutTemp       => PPCDMDCRDBUSOUT_OUT(30),
	Paths         => (0 => (CPMDCRCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCDMDCRDBUSOUT(31),
	GlitchData    => PPCDMDCRDBUSOUT31_GlitchData,
	OutSignalName => "PPCDMDCRDBUSOUT(31)",
	OutTemp       => PPCDMDCRDBUSOUT_OUT(31),
	Paths         => (0 => (CPMDCRCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCDMDCRREAD,
	GlitchData    => PPCDMDCRREAD_GlitchData,
	OutSignalName => "PPCDMDCRREAD",
	OutTemp       => PPCDMDCRREAD_OUT,
	Paths         => (0 => (CPMDCRCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCDMDCRUABUS(20),
	GlitchData    => PPCDMDCRUABUS20_GlitchData,
	OutSignalName => "PPCDMDCRUABUS(20)",
	OutTemp       => PPCDMDCRUABUS_OUT(20),
	Paths         => (0 => (CPMDCRCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCDMDCRUABUS(21),
	GlitchData    => PPCDMDCRUABUS21_GlitchData,
	OutSignalName => "PPCDMDCRUABUS(21)",
	OutTemp       => PPCDMDCRUABUS_OUT(21),
	Paths         => (0 => (CPMDCRCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCDMDCRWRITE,
	GlitchData    => PPCDMDCRWRITE_GlitchData,
	OutSignalName => "PPCDMDCRWRITE",
	OutTemp       => PPCDMDCRWRITE_OUT,
	Paths         => (0 => (CPMDCRCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCMPLBABORT,
	GlitchData    => PPCMPLBABORT_GlitchData,
	OutSignalName => "PPCMPLBABORT",
	OutTemp       => PPCMPLBABORT_OUT,
	Paths         => (0 => (CPMPPCMPLBCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCMPLBABUS(0),
	GlitchData    => PPCMPLBABUS0_GlitchData,
	OutSignalName => "PPCMPLBABUS(0)",
	OutTemp       => PPCMPLBABUS_OUT(0),
	Paths         => (0 => (CPMPPCMPLBCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCMPLBABUS(1),
	GlitchData    => PPCMPLBABUS1_GlitchData,
	OutSignalName => "PPCMPLBABUS(1)",
	OutTemp       => PPCMPLBABUS_OUT(1),
	Paths         => (0 => (CPMPPCMPLBCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCMPLBABUS(2),
	GlitchData    => PPCMPLBABUS2_GlitchData,
	OutSignalName => "PPCMPLBABUS(2)",
	OutTemp       => PPCMPLBABUS_OUT(2),
	Paths         => (0 => (CPMPPCMPLBCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCMPLBABUS(3),
	GlitchData    => PPCMPLBABUS3_GlitchData,
	OutSignalName => "PPCMPLBABUS(3)",
	OutTemp       => PPCMPLBABUS_OUT(3),
	Paths         => (0 => (CPMPPCMPLBCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCMPLBABUS(4),
	GlitchData    => PPCMPLBABUS4_GlitchData,
	OutSignalName => "PPCMPLBABUS(4)",
	OutTemp       => PPCMPLBABUS_OUT(4),
	Paths         => (0 => (CPMPPCMPLBCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCMPLBABUS(5),
	GlitchData    => PPCMPLBABUS5_GlitchData,
	OutSignalName => "PPCMPLBABUS(5)",
	OutTemp       => PPCMPLBABUS_OUT(5),
	Paths         => (0 => (CPMPPCMPLBCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCMPLBABUS(6),
	GlitchData    => PPCMPLBABUS6_GlitchData,
	OutSignalName => "PPCMPLBABUS(6)",
	OutTemp       => PPCMPLBABUS_OUT(6),
	Paths         => (0 => (CPMPPCMPLBCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCMPLBABUS(7),
	GlitchData    => PPCMPLBABUS7_GlitchData,
	OutSignalName => "PPCMPLBABUS(7)",
	OutTemp       => PPCMPLBABUS_OUT(7),
	Paths         => (0 => (CPMPPCMPLBCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCMPLBABUS(8),
	GlitchData    => PPCMPLBABUS8_GlitchData,
	OutSignalName => "PPCMPLBABUS(8)",
	OutTemp       => PPCMPLBABUS_OUT(8),
	Paths         => (0 => (CPMPPCMPLBCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCMPLBABUS(9),
	GlitchData    => PPCMPLBABUS9_GlitchData,
	OutSignalName => "PPCMPLBABUS(9)",
	OutTemp       => PPCMPLBABUS_OUT(9),
	Paths         => (0 => (CPMPPCMPLBCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCMPLBABUS(10),
	GlitchData    => PPCMPLBABUS10_GlitchData,
	OutSignalName => "PPCMPLBABUS(10)",
	OutTemp       => PPCMPLBABUS_OUT(10),
	Paths         => (0 => (CPMPPCMPLBCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCMPLBABUS(11),
	GlitchData    => PPCMPLBABUS11_GlitchData,
	OutSignalName => "PPCMPLBABUS(11)",
	OutTemp       => PPCMPLBABUS_OUT(11),
	Paths         => (0 => (CPMPPCMPLBCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCMPLBABUS(12),
	GlitchData    => PPCMPLBABUS12_GlitchData,
	OutSignalName => "PPCMPLBABUS(12)",
	OutTemp       => PPCMPLBABUS_OUT(12),
	Paths         => (0 => (CPMPPCMPLBCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCMPLBABUS(13),
	GlitchData    => PPCMPLBABUS13_GlitchData,
	OutSignalName => "PPCMPLBABUS(13)",
	OutTemp       => PPCMPLBABUS_OUT(13),
	Paths         => (0 => (CPMPPCMPLBCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCMPLBABUS(14),
	GlitchData    => PPCMPLBABUS14_GlitchData,
	OutSignalName => "PPCMPLBABUS(14)",
	OutTemp       => PPCMPLBABUS_OUT(14),
	Paths         => (0 => (CPMPPCMPLBCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCMPLBABUS(15),
	GlitchData    => PPCMPLBABUS15_GlitchData,
	OutSignalName => "PPCMPLBABUS(15)",
	OutTemp       => PPCMPLBABUS_OUT(15),
	Paths         => (0 => (CPMPPCMPLBCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCMPLBABUS(16),
	GlitchData    => PPCMPLBABUS16_GlitchData,
	OutSignalName => "PPCMPLBABUS(16)",
	OutTemp       => PPCMPLBABUS_OUT(16),
	Paths         => (0 => (CPMPPCMPLBCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCMPLBABUS(17),
	GlitchData    => PPCMPLBABUS17_GlitchData,
	OutSignalName => "PPCMPLBABUS(17)",
	OutTemp       => PPCMPLBABUS_OUT(17),
	Paths         => (0 => (CPMPPCMPLBCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCMPLBABUS(18),
	GlitchData    => PPCMPLBABUS18_GlitchData,
	OutSignalName => "PPCMPLBABUS(18)",
	OutTemp       => PPCMPLBABUS_OUT(18),
	Paths         => (0 => (CPMPPCMPLBCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCMPLBABUS(19),
	GlitchData    => PPCMPLBABUS19_GlitchData,
	OutSignalName => "PPCMPLBABUS(19)",
	OutTemp       => PPCMPLBABUS_OUT(19),
	Paths         => (0 => (CPMPPCMPLBCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCMPLBABUS(20),
	GlitchData    => PPCMPLBABUS20_GlitchData,
	OutSignalName => "PPCMPLBABUS(20)",
	OutTemp       => PPCMPLBABUS_OUT(20),
	Paths         => (0 => (CPMPPCMPLBCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCMPLBABUS(21),
	GlitchData    => PPCMPLBABUS21_GlitchData,
	OutSignalName => "PPCMPLBABUS(21)",
	OutTemp       => PPCMPLBABUS_OUT(21),
	Paths         => (0 => (CPMPPCMPLBCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCMPLBABUS(22),
	GlitchData    => PPCMPLBABUS22_GlitchData,
	OutSignalName => "PPCMPLBABUS(22)",
	OutTemp       => PPCMPLBABUS_OUT(22),
	Paths         => (0 => (CPMPPCMPLBCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCMPLBABUS(23),
	GlitchData    => PPCMPLBABUS23_GlitchData,
	OutSignalName => "PPCMPLBABUS(23)",
	OutTemp       => PPCMPLBABUS_OUT(23),
	Paths         => (0 => (CPMPPCMPLBCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCMPLBABUS(24),
	GlitchData    => PPCMPLBABUS24_GlitchData,
	OutSignalName => "PPCMPLBABUS(24)",
	OutTemp       => PPCMPLBABUS_OUT(24),
	Paths         => (0 => (CPMPPCMPLBCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCMPLBABUS(25),
	GlitchData    => PPCMPLBABUS25_GlitchData,
	OutSignalName => "PPCMPLBABUS(25)",
	OutTemp       => PPCMPLBABUS_OUT(25),
	Paths         => (0 => (CPMPPCMPLBCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCMPLBABUS(26),
	GlitchData    => PPCMPLBABUS26_GlitchData,
	OutSignalName => "PPCMPLBABUS(26)",
	OutTemp       => PPCMPLBABUS_OUT(26),
	Paths         => (0 => (CPMPPCMPLBCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCMPLBABUS(27),
	GlitchData    => PPCMPLBABUS27_GlitchData,
	OutSignalName => "PPCMPLBABUS(27)",
	OutTemp       => PPCMPLBABUS_OUT(27),
	Paths         => (0 => (CPMPPCMPLBCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCMPLBABUS(28),
	GlitchData    => PPCMPLBABUS28_GlitchData,
	OutSignalName => "PPCMPLBABUS(28)",
	OutTemp       => PPCMPLBABUS_OUT(28),
	Paths         => (0 => (CPMPPCMPLBCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCMPLBABUS(29),
	GlitchData    => PPCMPLBABUS29_GlitchData,
	OutSignalName => "PPCMPLBABUS(29)",
	OutTemp       => PPCMPLBABUS_OUT(29),
	Paths         => (0 => (CPMPPCMPLBCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCMPLBABUS(30),
	GlitchData    => PPCMPLBABUS30_GlitchData,
	OutSignalName => "PPCMPLBABUS(30)",
	OutTemp       => PPCMPLBABUS_OUT(30),
	Paths         => (0 => (CPMPPCMPLBCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCMPLBABUS(31),
	GlitchData    => PPCMPLBABUS31_GlitchData,
	OutSignalName => "PPCMPLBABUS(31)",
	OutTemp       => PPCMPLBABUS_OUT(31),
	Paths         => (0 => (CPMPPCMPLBCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCMPLBBE(0),
	GlitchData    => PPCMPLBBE0_GlitchData,
	OutSignalName => "PPCMPLBBE(0)",
	OutTemp       => PPCMPLBBE_OUT(0),
	Paths         => (0 => (CPMPPCMPLBCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCMPLBBE(1),
	GlitchData    => PPCMPLBBE1_GlitchData,
	OutSignalName => "PPCMPLBBE(1)",
	OutTemp       => PPCMPLBBE_OUT(1),
	Paths         => (0 => (CPMPPCMPLBCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCMPLBBE(2),
	GlitchData    => PPCMPLBBE2_GlitchData,
	OutSignalName => "PPCMPLBBE(2)",
	OutTemp       => PPCMPLBBE_OUT(2),
	Paths         => (0 => (CPMPPCMPLBCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCMPLBBE(3),
	GlitchData    => PPCMPLBBE3_GlitchData,
	OutSignalName => "PPCMPLBBE(3)",
	OutTemp       => PPCMPLBBE_OUT(3),
	Paths         => (0 => (CPMPPCMPLBCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCMPLBBE(4),
	GlitchData    => PPCMPLBBE4_GlitchData,
	OutSignalName => "PPCMPLBBE(4)",
	OutTemp       => PPCMPLBBE_OUT(4),
	Paths         => (0 => (CPMPPCMPLBCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCMPLBBE(5),
	GlitchData    => PPCMPLBBE5_GlitchData,
	OutSignalName => "PPCMPLBBE(5)",
	OutTemp       => PPCMPLBBE_OUT(5),
	Paths         => (0 => (CPMPPCMPLBCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCMPLBBE(6),
	GlitchData    => PPCMPLBBE6_GlitchData,
	OutSignalName => "PPCMPLBBE(6)",
	OutTemp       => PPCMPLBBE_OUT(6),
	Paths         => (0 => (CPMPPCMPLBCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCMPLBBE(7),
	GlitchData    => PPCMPLBBE7_GlitchData,
	OutSignalName => "PPCMPLBBE(7)",
	OutTemp       => PPCMPLBBE_OUT(7),
	Paths         => (0 => (CPMPPCMPLBCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCMPLBBE(8),
	GlitchData    => PPCMPLBBE8_GlitchData,
	OutSignalName => "PPCMPLBBE(8)",
	OutTemp       => PPCMPLBBE_OUT(8),
	Paths         => (0 => (CPMPPCMPLBCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCMPLBBE(9),
	GlitchData    => PPCMPLBBE9_GlitchData,
	OutSignalName => "PPCMPLBBE(9)",
	OutTemp       => PPCMPLBBE_OUT(9),
	Paths         => (0 => (CPMPPCMPLBCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCMPLBBE(10),
	GlitchData    => PPCMPLBBE10_GlitchData,
	OutSignalName => "PPCMPLBBE(10)",
	OutTemp       => PPCMPLBBE_OUT(10),
	Paths         => (0 => (CPMPPCMPLBCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCMPLBBE(11),
	GlitchData    => PPCMPLBBE11_GlitchData,
	OutSignalName => "PPCMPLBBE(11)",
	OutTemp       => PPCMPLBBE_OUT(11),
	Paths         => (0 => (CPMPPCMPLBCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCMPLBBE(12),
	GlitchData    => PPCMPLBBE12_GlitchData,
	OutSignalName => "PPCMPLBBE(12)",
	OutTemp       => PPCMPLBBE_OUT(12),
	Paths         => (0 => (CPMPPCMPLBCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCMPLBBE(13),
	GlitchData    => PPCMPLBBE13_GlitchData,
	OutSignalName => "PPCMPLBBE(13)",
	OutTemp       => PPCMPLBBE_OUT(13),
	Paths         => (0 => (CPMPPCMPLBCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCMPLBBE(14),
	GlitchData    => PPCMPLBBE14_GlitchData,
	OutSignalName => "PPCMPLBBE(14)",
	OutTemp       => PPCMPLBBE_OUT(14),
	Paths         => (0 => (CPMPPCMPLBCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCMPLBBE(15),
	GlitchData    => PPCMPLBBE15_GlitchData,
	OutSignalName => "PPCMPLBBE(15)",
	OutTemp       => PPCMPLBBE_OUT(15),
	Paths         => (0 => (CPMPPCMPLBCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCMPLBBUSLOCK,
	GlitchData    => PPCMPLBBUSLOCK_GlitchData,
	OutSignalName => "PPCMPLBBUSLOCK",
	OutTemp       => PPCMPLBBUSLOCK_OUT,
	Paths         => (0 => (CPMPPCMPLBCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCMPLBLOCKERR,
	GlitchData    => PPCMPLBLOCKERR_GlitchData,
	OutSignalName => "PPCMPLBLOCKERR",
	OutTemp       => PPCMPLBLOCKERR_OUT,
	Paths         => (0 => (CPMPPCMPLBCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCMPLBPRIORITY(0),
	GlitchData    => PPCMPLBPRIORITY0_GlitchData,
	OutSignalName => "PPCMPLBPRIORITY(0)",
	OutTemp       => PPCMPLBPRIORITY_OUT(0),
	Paths         => (0 => (CPMPPCMPLBCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCMPLBPRIORITY(1),
	GlitchData    => PPCMPLBPRIORITY1_GlitchData,
	OutSignalName => "PPCMPLBPRIORITY(1)",
	OutTemp       => PPCMPLBPRIORITY_OUT(1),
	Paths         => (0 => (CPMPPCMPLBCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCMPLBRDBURST,
	GlitchData    => PPCMPLBRDBURST_GlitchData,
	OutSignalName => "PPCMPLBRDBURST",
	OutTemp       => PPCMPLBRDBURST_OUT,
	Paths         => (0 => (CPMPPCMPLBCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCMPLBREQUEST,
	GlitchData    => PPCMPLBREQUEST_GlitchData,
	OutSignalName => "PPCMPLBREQUEST",
	OutTemp       => PPCMPLBREQUEST_OUT,
	Paths         => (0 => (CPMPPCMPLBCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCMPLBRNW,
	GlitchData    => PPCMPLBRNW_GlitchData,
	OutSignalName => "PPCMPLBRNW",
	OutTemp       => PPCMPLBRNW_OUT,
	Paths         => (0 => (CPMPPCMPLBCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCMPLBSIZE(0),
	GlitchData    => PPCMPLBSIZE0_GlitchData,
	OutSignalName => "PPCMPLBSIZE(0)",
	OutTemp       => PPCMPLBSIZE_OUT(0),
	Paths         => (0 => (CPMPPCMPLBCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCMPLBSIZE(1),
	GlitchData    => PPCMPLBSIZE1_GlitchData,
	OutSignalName => "PPCMPLBSIZE(1)",
	OutTemp       => PPCMPLBSIZE_OUT(1),
	Paths         => (0 => (CPMPPCMPLBCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCMPLBSIZE(2),
	GlitchData    => PPCMPLBSIZE2_GlitchData,
	OutSignalName => "PPCMPLBSIZE(2)",
	OutTemp       => PPCMPLBSIZE_OUT(2),
	Paths         => (0 => (CPMPPCMPLBCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCMPLBSIZE(3),
	GlitchData    => PPCMPLBSIZE3_GlitchData,
	OutSignalName => "PPCMPLBSIZE(3)",
	OutTemp       => PPCMPLBSIZE_OUT(3),
	Paths         => (0 => (CPMPPCMPLBCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCMPLBTATTRIBUTE(0),
	GlitchData    => PPCMPLBTATTRIBUTE0_GlitchData,
	OutSignalName => "PPCMPLBTATTRIBUTE(0)",
	OutTemp       => PPCMPLBTATTRIBUTE_OUT(0),
	Paths         => (0 => (CPMPPCMPLBCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCMPLBTATTRIBUTE(1),
	GlitchData    => PPCMPLBTATTRIBUTE1_GlitchData,
	OutSignalName => "PPCMPLBTATTRIBUTE(1)",
	OutTemp       => PPCMPLBTATTRIBUTE_OUT(1),
	Paths         => (0 => (CPMPPCMPLBCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCMPLBTATTRIBUTE(2),
	GlitchData    => PPCMPLBTATTRIBUTE2_GlitchData,
	OutSignalName => "PPCMPLBTATTRIBUTE(2)",
	OutTemp       => PPCMPLBTATTRIBUTE_OUT(2),
	Paths         => (0 => (CPMPPCMPLBCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCMPLBTATTRIBUTE(3),
	GlitchData    => PPCMPLBTATTRIBUTE3_GlitchData,
	OutSignalName => "PPCMPLBTATTRIBUTE(3)",
	OutTemp       => PPCMPLBTATTRIBUTE_OUT(3),
	Paths         => (0 => (CPMPPCMPLBCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCMPLBTATTRIBUTE(4),
	GlitchData    => PPCMPLBTATTRIBUTE4_GlitchData,
	OutSignalName => "PPCMPLBTATTRIBUTE(4)",
	OutTemp       => PPCMPLBTATTRIBUTE_OUT(4),
	Paths         => (0 => (CPMPPCMPLBCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCMPLBTATTRIBUTE(5),
	GlitchData    => PPCMPLBTATTRIBUTE5_GlitchData,
	OutSignalName => "PPCMPLBTATTRIBUTE(5)",
	OutTemp       => PPCMPLBTATTRIBUTE_OUT(5),
	Paths         => (0 => (CPMPPCMPLBCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCMPLBTATTRIBUTE(6),
	GlitchData    => PPCMPLBTATTRIBUTE6_GlitchData,
	OutSignalName => "PPCMPLBTATTRIBUTE(6)",
	OutTemp       => PPCMPLBTATTRIBUTE_OUT(6),
	Paths         => (0 => (CPMPPCMPLBCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCMPLBTATTRIBUTE(7),
	GlitchData    => PPCMPLBTATTRIBUTE7_GlitchData,
	OutSignalName => "PPCMPLBTATTRIBUTE(7)",
	OutTemp       => PPCMPLBTATTRIBUTE_OUT(7),
	Paths         => (0 => (CPMPPCMPLBCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCMPLBTATTRIBUTE(8),
	GlitchData    => PPCMPLBTATTRIBUTE8_GlitchData,
	OutSignalName => "PPCMPLBTATTRIBUTE(8)",
	OutTemp       => PPCMPLBTATTRIBUTE_OUT(8),
	Paths         => (0 => (CPMPPCMPLBCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCMPLBTATTRIBUTE(9),
	GlitchData    => PPCMPLBTATTRIBUTE9_GlitchData,
	OutSignalName => "PPCMPLBTATTRIBUTE(9)",
	OutTemp       => PPCMPLBTATTRIBUTE_OUT(9),
	Paths         => (0 => (CPMPPCMPLBCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCMPLBTATTRIBUTE(10),
	GlitchData    => PPCMPLBTATTRIBUTE10_GlitchData,
	OutSignalName => "PPCMPLBTATTRIBUTE(10)",
	OutTemp       => PPCMPLBTATTRIBUTE_OUT(10),
	Paths         => (0 => (CPMPPCMPLBCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCMPLBTATTRIBUTE(11),
	GlitchData    => PPCMPLBTATTRIBUTE11_GlitchData,
	OutSignalName => "PPCMPLBTATTRIBUTE(11)",
	OutTemp       => PPCMPLBTATTRIBUTE_OUT(11),
	Paths         => (0 => (CPMPPCMPLBCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCMPLBTATTRIBUTE(12),
	GlitchData    => PPCMPLBTATTRIBUTE12_GlitchData,
	OutSignalName => "PPCMPLBTATTRIBUTE(12)",
	OutTemp       => PPCMPLBTATTRIBUTE_OUT(12),
	Paths         => (0 => (CPMPPCMPLBCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCMPLBTATTRIBUTE(13),
	GlitchData    => PPCMPLBTATTRIBUTE13_GlitchData,
	OutSignalName => "PPCMPLBTATTRIBUTE(13)",
	OutTemp       => PPCMPLBTATTRIBUTE_OUT(13),
	Paths         => (0 => (CPMPPCMPLBCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCMPLBTATTRIBUTE(14),
	GlitchData    => PPCMPLBTATTRIBUTE14_GlitchData,
	OutSignalName => "PPCMPLBTATTRIBUTE(14)",
	OutTemp       => PPCMPLBTATTRIBUTE_OUT(14),
	Paths         => (0 => (CPMPPCMPLBCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCMPLBTATTRIBUTE(15),
	GlitchData    => PPCMPLBTATTRIBUTE15_GlitchData,
	OutSignalName => "PPCMPLBTATTRIBUTE(15)",
	OutTemp       => PPCMPLBTATTRIBUTE_OUT(15),
	Paths         => (0 => (CPMPPCMPLBCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCMPLBTYPE(0),
	GlitchData    => PPCMPLBTYPE0_GlitchData,
	OutSignalName => "PPCMPLBTYPE(0)",
	OutTemp       => PPCMPLBTYPE_OUT(0),
	Paths         => (0 => (CPMPPCMPLBCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCMPLBTYPE(1),
	GlitchData    => PPCMPLBTYPE1_GlitchData,
	OutSignalName => "PPCMPLBTYPE(1)",
	OutTemp       => PPCMPLBTYPE_OUT(1),
	Paths         => (0 => (CPMPPCMPLBCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCMPLBTYPE(2),
	GlitchData    => PPCMPLBTYPE2_GlitchData,
	OutSignalName => "PPCMPLBTYPE(2)",
	OutTemp       => PPCMPLBTYPE_OUT(2),
	Paths         => (0 => (CPMPPCMPLBCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCMPLBUABUS(28),
	GlitchData    => PPCMPLBUABUS28_GlitchData,
	OutSignalName => "PPCMPLBUABUS(28)",
	OutTemp       => PPCMPLBUABUS_OUT(28),
	Paths         => (0 => (CPMPPCMPLBCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCMPLBUABUS(29),
	GlitchData    => PPCMPLBUABUS29_GlitchData,
	OutSignalName => "PPCMPLBUABUS(29)",
	OutTemp       => PPCMPLBUABUS_OUT(29),
	Paths         => (0 => (CPMPPCMPLBCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCMPLBUABUS(30),
	GlitchData    => PPCMPLBUABUS30_GlitchData,
	OutSignalName => "PPCMPLBUABUS(30)",
	OutTemp       => PPCMPLBUABUS_OUT(30),
	Paths         => (0 => (CPMPPCMPLBCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCMPLBUABUS(31),
	GlitchData    => PPCMPLBUABUS31_GlitchData,
	OutSignalName => "PPCMPLBUABUS(31)",
	OutTemp       => PPCMPLBUABUS_OUT(31),
	Paths         => (0 => (CPMPPCMPLBCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCMPLBWRBURST,
	GlitchData    => PPCMPLBWRBURST_GlitchData,
	OutSignalName => "PPCMPLBWRBURST",
	OutTemp       => PPCMPLBWRBURST_OUT,
	Paths         => (0 => (CPMPPCMPLBCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCMPLBWRDBUS(0),
	GlitchData    => PPCMPLBWRDBUS0_GlitchData,
	OutSignalName => "PPCMPLBWRDBUS(0)",
	OutTemp       => PPCMPLBWRDBUS_OUT(0),
	Paths         => (0 => (CPMPPCMPLBCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCMPLBWRDBUS(1),
	GlitchData    => PPCMPLBWRDBUS1_GlitchData,
	OutSignalName => "PPCMPLBWRDBUS(1)",
	OutTemp       => PPCMPLBWRDBUS_OUT(1),
	Paths         => (0 => (CPMPPCMPLBCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCMPLBWRDBUS(2),
	GlitchData    => PPCMPLBWRDBUS2_GlitchData,
	OutSignalName => "PPCMPLBWRDBUS(2)",
	OutTemp       => PPCMPLBWRDBUS_OUT(2),
	Paths         => (0 => (CPMPPCMPLBCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCMPLBWRDBUS(3),
	GlitchData    => PPCMPLBWRDBUS3_GlitchData,
	OutSignalName => "PPCMPLBWRDBUS(3)",
	OutTemp       => PPCMPLBWRDBUS_OUT(3),
	Paths         => (0 => (CPMPPCMPLBCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCMPLBWRDBUS(4),
	GlitchData    => PPCMPLBWRDBUS4_GlitchData,
	OutSignalName => "PPCMPLBWRDBUS(4)",
	OutTemp       => PPCMPLBWRDBUS_OUT(4),
	Paths         => (0 => (CPMPPCMPLBCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCMPLBWRDBUS(5),
	GlitchData    => PPCMPLBWRDBUS5_GlitchData,
	OutSignalName => "PPCMPLBWRDBUS(5)",
	OutTemp       => PPCMPLBWRDBUS_OUT(5),
	Paths         => (0 => (CPMPPCMPLBCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCMPLBWRDBUS(6),
	GlitchData    => PPCMPLBWRDBUS6_GlitchData,
	OutSignalName => "PPCMPLBWRDBUS(6)",
	OutTemp       => PPCMPLBWRDBUS_OUT(6),
	Paths         => (0 => (CPMPPCMPLBCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCMPLBWRDBUS(7),
	GlitchData    => PPCMPLBWRDBUS7_GlitchData,
	OutSignalName => "PPCMPLBWRDBUS(7)",
	OutTemp       => PPCMPLBWRDBUS_OUT(7),
	Paths         => (0 => (CPMPPCMPLBCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCMPLBWRDBUS(8),
	GlitchData    => PPCMPLBWRDBUS8_GlitchData,
	OutSignalName => "PPCMPLBWRDBUS(8)",
	OutTemp       => PPCMPLBWRDBUS_OUT(8),
	Paths         => (0 => (CPMPPCMPLBCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCMPLBWRDBUS(9),
	GlitchData    => PPCMPLBWRDBUS9_GlitchData,
	OutSignalName => "PPCMPLBWRDBUS(9)",
	OutTemp       => PPCMPLBWRDBUS_OUT(9),
	Paths         => (0 => (CPMPPCMPLBCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCMPLBWRDBUS(10),
	GlitchData    => PPCMPLBWRDBUS10_GlitchData,
	OutSignalName => "PPCMPLBWRDBUS(10)",
	OutTemp       => PPCMPLBWRDBUS_OUT(10),
	Paths         => (0 => (CPMPPCMPLBCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCMPLBWRDBUS(11),
	GlitchData    => PPCMPLBWRDBUS11_GlitchData,
	OutSignalName => "PPCMPLBWRDBUS(11)",
	OutTemp       => PPCMPLBWRDBUS_OUT(11),
	Paths         => (0 => (CPMPPCMPLBCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCMPLBWRDBUS(12),
	GlitchData    => PPCMPLBWRDBUS12_GlitchData,
	OutSignalName => "PPCMPLBWRDBUS(12)",
	OutTemp       => PPCMPLBWRDBUS_OUT(12),
	Paths         => (0 => (CPMPPCMPLBCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCMPLBWRDBUS(13),
	GlitchData    => PPCMPLBWRDBUS13_GlitchData,
	OutSignalName => "PPCMPLBWRDBUS(13)",
	OutTemp       => PPCMPLBWRDBUS_OUT(13),
	Paths         => (0 => (CPMPPCMPLBCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCMPLBWRDBUS(14),
	GlitchData    => PPCMPLBWRDBUS14_GlitchData,
	OutSignalName => "PPCMPLBWRDBUS(14)",
	OutTemp       => PPCMPLBWRDBUS_OUT(14),
	Paths         => (0 => (CPMPPCMPLBCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCMPLBWRDBUS(15),
	GlitchData    => PPCMPLBWRDBUS15_GlitchData,
	OutSignalName => "PPCMPLBWRDBUS(15)",
	OutTemp       => PPCMPLBWRDBUS_OUT(15),
	Paths         => (0 => (CPMPPCMPLBCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCMPLBWRDBUS(16),
	GlitchData    => PPCMPLBWRDBUS16_GlitchData,
	OutSignalName => "PPCMPLBWRDBUS(16)",
	OutTemp       => PPCMPLBWRDBUS_OUT(16),
	Paths         => (0 => (CPMPPCMPLBCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCMPLBWRDBUS(17),
	GlitchData    => PPCMPLBWRDBUS17_GlitchData,
	OutSignalName => "PPCMPLBWRDBUS(17)",
	OutTemp       => PPCMPLBWRDBUS_OUT(17),
	Paths         => (0 => (CPMPPCMPLBCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCMPLBWRDBUS(18),
	GlitchData    => PPCMPLBWRDBUS18_GlitchData,
	OutSignalName => "PPCMPLBWRDBUS(18)",
	OutTemp       => PPCMPLBWRDBUS_OUT(18),
	Paths         => (0 => (CPMPPCMPLBCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCMPLBWRDBUS(19),
	GlitchData    => PPCMPLBWRDBUS19_GlitchData,
	OutSignalName => "PPCMPLBWRDBUS(19)",
	OutTemp       => PPCMPLBWRDBUS_OUT(19),
	Paths         => (0 => (CPMPPCMPLBCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCMPLBWRDBUS(20),
	GlitchData    => PPCMPLBWRDBUS20_GlitchData,
	OutSignalName => "PPCMPLBWRDBUS(20)",
	OutTemp       => PPCMPLBWRDBUS_OUT(20),
	Paths         => (0 => (CPMPPCMPLBCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCMPLBWRDBUS(21),
	GlitchData    => PPCMPLBWRDBUS21_GlitchData,
	OutSignalName => "PPCMPLBWRDBUS(21)",
	OutTemp       => PPCMPLBWRDBUS_OUT(21),
	Paths         => (0 => (CPMPPCMPLBCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCMPLBWRDBUS(22),
	GlitchData    => PPCMPLBWRDBUS22_GlitchData,
	OutSignalName => "PPCMPLBWRDBUS(22)",
	OutTemp       => PPCMPLBWRDBUS_OUT(22),
	Paths         => (0 => (CPMPPCMPLBCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCMPLBWRDBUS(23),
	GlitchData    => PPCMPLBWRDBUS23_GlitchData,
	OutSignalName => "PPCMPLBWRDBUS(23)",
	OutTemp       => PPCMPLBWRDBUS_OUT(23),
	Paths         => (0 => (CPMPPCMPLBCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCMPLBWRDBUS(24),
	GlitchData    => PPCMPLBWRDBUS24_GlitchData,
	OutSignalName => "PPCMPLBWRDBUS(24)",
	OutTemp       => PPCMPLBWRDBUS_OUT(24),
	Paths         => (0 => (CPMPPCMPLBCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCMPLBWRDBUS(25),
	GlitchData    => PPCMPLBWRDBUS25_GlitchData,
	OutSignalName => "PPCMPLBWRDBUS(25)",
	OutTemp       => PPCMPLBWRDBUS_OUT(25),
	Paths         => (0 => (CPMPPCMPLBCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCMPLBWRDBUS(26),
	GlitchData    => PPCMPLBWRDBUS26_GlitchData,
	OutSignalName => "PPCMPLBWRDBUS(26)",
	OutTemp       => PPCMPLBWRDBUS_OUT(26),
	Paths         => (0 => (CPMPPCMPLBCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCMPLBWRDBUS(27),
	GlitchData    => PPCMPLBWRDBUS27_GlitchData,
	OutSignalName => "PPCMPLBWRDBUS(27)",
	OutTemp       => PPCMPLBWRDBUS_OUT(27),
	Paths         => (0 => (CPMPPCMPLBCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCMPLBWRDBUS(28),
	GlitchData    => PPCMPLBWRDBUS28_GlitchData,
	OutSignalName => "PPCMPLBWRDBUS(28)",
	OutTemp       => PPCMPLBWRDBUS_OUT(28),
	Paths         => (0 => (CPMPPCMPLBCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCMPLBWRDBUS(29),
	GlitchData    => PPCMPLBWRDBUS29_GlitchData,
	OutSignalName => "PPCMPLBWRDBUS(29)",
	OutTemp       => PPCMPLBWRDBUS_OUT(29),
	Paths         => (0 => (CPMPPCMPLBCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCMPLBWRDBUS(30),
	GlitchData    => PPCMPLBWRDBUS30_GlitchData,
	OutSignalName => "PPCMPLBWRDBUS(30)",
	OutTemp       => PPCMPLBWRDBUS_OUT(30),
	Paths         => (0 => (CPMPPCMPLBCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCMPLBWRDBUS(31),
	GlitchData    => PPCMPLBWRDBUS31_GlitchData,
	OutSignalName => "PPCMPLBWRDBUS(31)",
	OutTemp       => PPCMPLBWRDBUS_OUT(31),
	Paths         => (0 => (CPMPPCMPLBCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCMPLBWRDBUS(32),
	GlitchData    => PPCMPLBWRDBUS32_GlitchData,
	OutSignalName => "PPCMPLBWRDBUS(32)",
	OutTemp       => PPCMPLBWRDBUS_OUT(32),
	Paths         => (0 => (CPMPPCMPLBCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCMPLBWRDBUS(33),
	GlitchData    => PPCMPLBWRDBUS33_GlitchData,
	OutSignalName => "PPCMPLBWRDBUS(33)",
	OutTemp       => PPCMPLBWRDBUS_OUT(33),
	Paths         => (0 => (CPMPPCMPLBCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCMPLBWRDBUS(34),
	GlitchData    => PPCMPLBWRDBUS34_GlitchData,
	OutSignalName => "PPCMPLBWRDBUS(34)",
	OutTemp       => PPCMPLBWRDBUS_OUT(34),
	Paths         => (0 => (CPMPPCMPLBCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCMPLBWRDBUS(35),
	GlitchData    => PPCMPLBWRDBUS35_GlitchData,
	OutSignalName => "PPCMPLBWRDBUS(35)",
	OutTemp       => PPCMPLBWRDBUS_OUT(35),
	Paths         => (0 => (CPMPPCMPLBCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCMPLBWRDBUS(36),
	GlitchData    => PPCMPLBWRDBUS36_GlitchData,
	OutSignalName => "PPCMPLBWRDBUS(36)",
	OutTemp       => PPCMPLBWRDBUS_OUT(36),
	Paths         => (0 => (CPMPPCMPLBCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCMPLBWRDBUS(37),
	GlitchData    => PPCMPLBWRDBUS37_GlitchData,
	OutSignalName => "PPCMPLBWRDBUS(37)",
	OutTemp       => PPCMPLBWRDBUS_OUT(37),
	Paths         => (0 => (CPMPPCMPLBCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCMPLBWRDBUS(38),
	GlitchData    => PPCMPLBWRDBUS38_GlitchData,
	OutSignalName => "PPCMPLBWRDBUS(38)",
	OutTemp       => PPCMPLBWRDBUS_OUT(38),
	Paths         => (0 => (CPMPPCMPLBCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCMPLBWRDBUS(39),
	GlitchData    => PPCMPLBWRDBUS39_GlitchData,
	OutSignalName => "PPCMPLBWRDBUS(39)",
	OutTemp       => PPCMPLBWRDBUS_OUT(39),
	Paths         => (0 => (CPMPPCMPLBCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCMPLBWRDBUS(40),
	GlitchData    => PPCMPLBWRDBUS40_GlitchData,
	OutSignalName => "PPCMPLBWRDBUS(40)",
	OutTemp       => PPCMPLBWRDBUS_OUT(40),
	Paths         => (0 => (CPMPPCMPLBCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCMPLBWRDBUS(41),
	GlitchData    => PPCMPLBWRDBUS41_GlitchData,
	OutSignalName => "PPCMPLBWRDBUS(41)",
	OutTemp       => PPCMPLBWRDBUS_OUT(41),
	Paths         => (0 => (CPMPPCMPLBCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCMPLBWRDBUS(42),
	GlitchData    => PPCMPLBWRDBUS42_GlitchData,
	OutSignalName => "PPCMPLBWRDBUS(42)",
	OutTemp       => PPCMPLBWRDBUS_OUT(42),
	Paths         => (0 => (CPMPPCMPLBCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCMPLBWRDBUS(43),
	GlitchData    => PPCMPLBWRDBUS43_GlitchData,
	OutSignalName => "PPCMPLBWRDBUS(43)",
	OutTemp       => PPCMPLBWRDBUS_OUT(43),
	Paths         => (0 => (CPMPPCMPLBCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCMPLBWRDBUS(44),
	GlitchData    => PPCMPLBWRDBUS44_GlitchData,
	OutSignalName => "PPCMPLBWRDBUS(44)",
	OutTemp       => PPCMPLBWRDBUS_OUT(44),
	Paths         => (0 => (CPMPPCMPLBCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCMPLBWRDBUS(45),
	GlitchData    => PPCMPLBWRDBUS45_GlitchData,
	OutSignalName => "PPCMPLBWRDBUS(45)",
	OutTemp       => PPCMPLBWRDBUS_OUT(45),
	Paths         => (0 => (CPMPPCMPLBCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCMPLBWRDBUS(46),
	GlitchData    => PPCMPLBWRDBUS46_GlitchData,
	OutSignalName => "PPCMPLBWRDBUS(46)",
	OutTemp       => PPCMPLBWRDBUS_OUT(46),
	Paths         => (0 => (CPMPPCMPLBCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCMPLBWRDBUS(47),
	GlitchData    => PPCMPLBWRDBUS47_GlitchData,
	OutSignalName => "PPCMPLBWRDBUS(47)",
	OutTemp       => PPCMPLBWRDBUS_OUT(47),
	Paths         => (0 => (CPMPPCMPLBCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCMPLBWRDBUS(48),
	GlitchData    => PPCMPLBWRDBUS48_GlitchData,
	OutSignalName => "PPCMPLBWRDBUS(48)",
	OutTemp       => PPCMPLBWRDBUS_OUT(48),
	Paths         => (0 => (CPMPPCMPLBCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCMPLBWRDBUS(49),
	GlitchData    => PPCMPLBWRDBUS49_GlitchData,
	OutSignalName => "PPCMPLBWRDBUS(49)",
	OutTemp       => PPCMPLBWRDBUS_OUT(49),
	Paths         => (0 => (CPMPPCMPLBCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCMPLBWRDBUS(50),
	GlitchData    => PPCMPLBWRDBUS50_GlitchData,
	OutSignalName => "PPCMPLBWRDBUS(50)",
	OutTemp       => PPCMPLBWRDBUS_OUT(50),
	Paths         => (0 => (CPMPPCMPLBCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCMPLBWRDBUS(51),
	GlitchData    => PPCMPLBWRDBUS51_GlitchData,
	OutSignalName => "PPCMPLBWRDBUS(51)",
	OutTemp       => PPCMPLBWRDBUS_OUT(51),
	Paths         => (0 => (CPMPPCMPLBCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCMPLBWRDBUS(52),
	GlitchData    => PPCMPLBWRDBUS52_GlitchData,
	OutSignalName => "PPCMPLBWRDBUS(52)",
	OutTemp       => PPCMPLBWRDBUS_OUT(52),
	Paths         => (0 => (CPMPPCMPLBCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCMPLBWRDBUS(53),
	GlitchData    => PPCMPLBWRDBUS53_GlitchData,
	OutSignalName => "PPCMPLBWRDBUS(53)",
	OutTemp       => PPCMPLBWRDBUS_OUT(53),
	Paths         => (0 => (CPMPPCMPLBCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCMPLBWRDBUS(54),
	GlitchData    => PPCMPLBWRDBUS54_GlitchData,
	OutSignalName => "PPCMPLBWRDBUS(54)",
	OutTemp       => PPCMPLBWRDBUS_OUT(54),
	Paths         => (0 => (CPMPPCMPLBCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCMPLBWRDBUS(55),
	GlitchData    => PPCMPLBWRDBUS55_GlitchData,
	OutSignalName => "PPCMPLBWRDBUS(55)",
	OutTemp       => PPCMPLBWRDBUS_OUT(55),
	Paths         => (0 => (CPMPPCMPLBCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCMPLBWRDBUS(56),
	GlitchData    => PPCMPLBWRDBUS56_GlitchData,
	OutSignalName => "PPCMPLBWRDBUS(56)",
	OutTemp       => PPCMPLBWRDBUS_OUT(56),
	Paths         => (0 => (CPMPPCMPLBCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCMPLBWRDBUS(57),
	GlitchData    => PPCMPLBWRDBUS57_GlitchData,
	OutSignalName => "PPCMPLBWRDBUS(57)",
	OutTemp       => PPCMPLBWRDBUS_OUT(57),
	Paths         => (0 => (CPMPPCMPLBCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCMPLBWRDBUS(58),
	GlitchData    => PPCMPLBWRDBUS58_GlitchData,
	OutSignalName => "PPCMPLBWRDBUS(58)",
	OutTemp       => PPCMPLBWRDBUS_OUT(58),
	Paths         => (0 => (CPMPPCMPLBCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCMPLBWRDBUS(59),
	GlitchData    => PPCMPLBWRDBUS59_GlitchData,
	OutSignalName => "PPCMPLBWRDBUS(59)",
	OutTemp       => PPCMPLBWRDBUS_OUT(59),
	Paths         => (0 => (CPMPPCMPLBCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCMPLBWRDBUS(60),
	GlitchData    => PPCMPLBWRDBUS60_GlitchData,
	OutSignalName => "PPCMPLBWRDBUS(60)",
	OutTemp       => PPCMPLBWRDBUS_OUT(60),
	Paths         => (0 => (CPMPPCMPLBCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCMPLBWRDBUS(61),
	GlitchData    => PPCMPLBWRDBUS61_GlitchData,
	OutSignalName => "PPCMPLBWRDBUS(61)",
	OutTemp       => PPCMPLBWRDBUS_OUT(61),
	Paths         => (0 => (CPMPPCMPLBCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCMPLBWRDBUS(62),
	GlitchData    => PPCMPLBWRDBUS62_GlitchData,
	OutSignalName => "PPCMPLBWRDBUS(62)",
	OutTemp       => PPCMPLBWRDBUS_OUT(62),
	Paths         => (0 => (CPMPPCMPLBCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCMPLBWRDBUS(63),
	GlitchData    => PPCMPLBWRDBUS63_GlitchData,
	OutSignalName => "PPCMPLBWRDBUS(63)",
	OutTemp       => PPCMPLBWRDBUS_OUT(63),
	Paths         => (0 => (CPMPPCMPLBCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCMPLBWRDBUS(64),
	GlitchData    => PPCMPLBWRDBUS64_GlitchData,
	OutSignalName => "PPCMPLBWRDBUS(64)",
	OutTemp       => PPCMPLBWRDBUS_OUT(64),
	Paths         => (0 => (CPMPPCMPLBCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCMPLBWRDBUS(65),
	GlitchData    => PPCMPLBWRDBUS65_GlitchData,
	OutSignalName => "PPCMPLBWRDBUS(65)",
	OutTemp       => PPCMPLBWRDBUS_OUT(65),
	Paths         => (0 => (CPMPPCMPLBCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCMPLBWRDBUS(66),
	GlitchData    => PPCMPLBWRDBUS66_GlitchData,
	OutSignalName => "PPCMPLBWRDBUS(66)",
	OutTemp       => PPCMPLBWRDBUS_OUT(66),
	Paths         => (0 => (CPMPPCMPLBCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCMPLBWRDBUS(67),
	GlitchData    => PPCMPLBWRDBUS67_GlitchData,
	OutSignalName => "PPCMPLBWRDBUS(67)",
	OutTemp       => PPCMPLBWRDBUS_OUT(67),
	Paths         => (0 => (CPMPPCMPLBCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCMPLBWRDBUS(68),
	GlitchData    => PPCMPLBWRDBUS68_GlitchData,
	OutSignalName => "PPCMPLBWRDBUS(68)",
	OutTemp       => PPCMPLBWRDBUS_OUT(68),
	Paths         => (0 => (CPMPPCMPLBCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCMPLBWRDBUS(69),
	GlitchData    => PPCMPLBWRDBUS69_GlitchData,
	OutSignalName => "PPCMPLBWRDBUS(69)",
	OutTemp       => PPCMPLBWRDBUS_OUT(69),
	Paths         => (0 => (CPMPPCMPLBCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCMPLBWRDBUS(70),
	GlitchData    => PPCMPLBWRDBUS70_GlitchData,
	OutSignalName => "PPCMPLBWRDBUS(70)",
	OutTemp       => PPCMPLBWRDBUS_OUT(70),
	Paths         => (0 => (CPMPPCMPLBCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCMPLBWRDBUS(71),
	GlitchData    => PPCMPLBWRDBUS71_GlitchData,
	OutSignalName => "PPCMPLBWRDBUS(71)",
	OutTemp       => PPCMPLBWRDBUS_OUT(71),
	Paths         => (0 => (CPMPPCMPLBCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCMPLBWRDBUS(72),
	GlitchData    => PPCMPLBWRDBUS72_GlitchData,
	OutSignalName => "PPCMPLBWRDBUS(72)",
	OutTemp       => PPCMPLBWRDBUS_OUT(72),
	Paths         => (0 => (CPMPPCMPLBCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCMPLBWRDBUS(73),
	GlitchData    => PPCMPLBWRDBUS73_GlitchData,
	OutSignalName => "PPCMPLBWRDBUS(73)",
	OutTemp       => PPCMPLBWRDBUS_OUT(73),
	Paths         => (0 => (CPMPPCMPLBCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCMPLBWRDBUS(74),
	GlitchData    => PPCMPLBWRDBUS74_GlitchData,
	OutSignalName => "PPCMPLBWRDBUS(74)",
	OutTemp       => PPCMPLBWRDBUS_OUT(74),
	Paths         => (0 => (CPMPPCMPLBCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCMPLBWRDBUS(75),
	GlitchData    => PPCMPLBWRDBUS75_GlitchData,
	OutSignalName => "PPCMPLBWRDBUS(75)",
	OutTemp       => PPCMPLBWRDBUS_OUT(75),
	Paths         => (0 => (CPMPPCMPLBCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCMPLBWRDBUS(76),
	GlitchData    => PPCMPLBWRDBUS76_GlitchData,
	OutSignalName => "PPCMPLBWRDBUS(76)",
	OutTemp       => PPCMPLBWRDBUS_OUT(76),
	Paths         => (0 => (CPMPPCMPLBCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCMPLBWRDBUS(77),
	GlitchData    => PPCMPLBWRDBUS77_GlitchData,
	OutSignalName => "PPCMPLBWRDBUS(77)",
	OutTemp       => PPCMPLBWRDBUS_OUT(77),
	Paths         => (0 => (CPMPPCMPLBCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCMPLBWRDBUS(78),
	GlitchData    => PPCMPLBWRDBUS78_GlitchData,
	OutSignalName => "PPCMPLBWRDBUS(78)",
	OutTemp       => PPCMPLBWRDBUS_OUT(78),
	Paths         => (0 => (CPMPPCMPLBCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCMPLBWRDBUS(79),
	GlitchData    => PPCMPLBWRDBUS79_GlitchData,
	OutSignalName => "PPCMPLBWRDBUS(79)",
	OutTemp       => PPCMPLBWRDBUS_OUT(79),
	Paths         => (0 => (CPMPPCMPLBCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCMPLBWRDBUS(80),
	GlitchData    => PPCMPLBWRDBUS80_GlitchData,
	OutSignalName => "PPCMPLBWRDBUS(80)",
	OutTemp       => PPCMPLBWRDBUS_OUT(80),
	Paths         => (0 => (CPMPPCMPLBCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCMPLBWRDBUS(81),
	GlitchData    => PPCMPLBWRDBUS81_GlitchData,
	OutSignalName => "PPCMPLBWRDBUS(81)",
	OutTemp       => PPCMPLBWRDBUS_OUT(81),
	Paths         => (0 => (CPMPPCMPLBCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCMPLBWRDBUS(82),
	GlitchData    => PPCMPLBWRDBUS82_GlitchData,
	OutSignalName => "PPCMPLBWRDBUS(82)",
	OutTemp       => PPCMPLBWRDBUS_OUT(82),
	Paths         => (0 => (CPMPPCMPLBCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCMPLBWRDBUS(83),
	GlitchData    => PPCMPLBWRDBUS83_GlitchData,
	OutSignalName => "PPCMPLBWRDBUS(83)",
	OutTemp       => PPCMPLBWRDBUS_OUT(83),
	Paths         => (0 => (CPMPPCMPLBCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCMPLBWRDBUS(84),
	GlitchData    => PPCMPLBWRDBUS84_GlitchData,
	OutSignalName => "PPCMPLBWRDBUS(84)",
	OutTemp       => PPCMPLBWRDBUS_OUT(84),
	Paths         => (0 => (CPMPPCMPLBCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCMPLBWRDBUS(85),
	GlitchData    => PPCMPLBWRDBUS85_GlitchData,
	OutSignalName => "PPCMPLBWRDBUS(85)",
	OutTemp       => PPCMPLBWRDBUS_OUT(85),
	Paths         => (0 => (CPMPPCMPLBCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCMPLBWRDBUS(86),
	GlitchData    => PPCMPLBWRDBUS86_GlitchData,
	OutSignalName => "PPCMPLBWRDBUS(86)",
	OutTemp       => PPCMPLBWRDBUS_OUT(86),
	Paths         => (0 => (CPMPPCMPLBCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCMPLBWRDBUS(87),
	GlitchData    => PPCMPLBWRDBUS87_GlitchData,
	OutSignalName => "PPCMPLBWRDBUS(87)",
	OutTemp       => PPCMPLBWRDBUS_OUT(87),
	Paths         => (0 => (CPMPPCMPLBCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCMPLBWRDBUS(88),
	GlitchData    => PPCMPLBWRDBUS88_GlitchData,
	OutSignalName => "PPCMPLBWRDBUS(88)",
	OutTemp       => PPCMPLBWRDBUS_OUT(88),
	Paths         => (0 => (CPMPPCMPLBCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCMPLBWRDBUS(89),
	GlitchData    => PPCMPLBWRDBUS89_GlitchData,
	OutSignalName => "PPCMPLBWRDBUS(89)",
	OutTemp       => PPCMPLBWRDBUS_OUT(89),
	Paths         => (0 => (CPMPPCMPLBCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCMPLBWRDBUS(90),
	GlitchData    => PPCMPLBWRDBUS90_GlitchData,
	OutSignalName => "PPCMPLBWRDBUS(90)",
	OutTemp       => PPCMPLBWRDBUS_OUT(90),
	Paths         => (0 => (CPMPPCMPLBCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCMPLBWRDBUS(91),
	GlitchData    => PPCMPLBWRDBUS91_GlitchData,
	OutSignalName => "PPCMPLBWRDBUS(91)",
	OutTemp       => PPCMPLBWRDBUS_OUT(91),
	Paths         => (0 => (CPMPPCMPLBCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCMPLBWRDBUS(92),
	GlitchData    => PPCMPLBWRDBUS92_GlitchData,
	OutSignalName => "PPCMPLBWRDBUS(92)",
	OutTemp       => PPCMPLBWRDBUS_OUT(92),
	Paths         => (0 => (CPMPPCMPLBCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCMPLBWRDBUS(93),
	GlitchData    => PPCMPLBWRDBUS93_GlitchData,
	OutSignalName => "PPCMPLBWRDBUS(93)",
	OutTemp       => PPCMPLBWRDBUS_OUT(93),
	Paths         => (0 => (CPMPPCMPLBCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCMPLBWRDBUS(94),
	GlitchData    => PPCMPLBWRDBUS94_GlitchData,
	OutSignalName => "PPCMPLBWRDBUS(94)",
	OutTemp       => PPCMPLBWRDBUS_OUT(94),
	Paths         => (0 => (CPMPPCMPLBCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCMPLBWRDBUS(95),
	GlitchData    => PPCMPLBWRDBUS95_GlitchData,
	OutSignalName => "PPCMPLBWRDBUS(95)",
	OutTemp       => PPCMPLBWRDBUS_OUT(95),
	Paths         => (0 => (CPMPPCMPLBCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCMPLBWRDBUS(96),
	GlitchData    => PPCMPLBWRDBUS96_GlitchData,
	OutSignalName => "PPCMPLBWRDBUS(96)",
	OutTemp       => PPCMPLBWRDBUS_OUT(96),
	Paths         => (0 => (CPMPPCMPLBCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCMPLBWRDBUS(97),
	GlitchData    => PPCMPLBWRDBUS97_GlitchData,
	OutSignalName => "PPCMPLBWRDBUS(97)",
	OutTemp       => PPCMPLBWRDBUS_OUT(97),
	Paths         => (0 => (CPMPPCMPLBCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCMPLBWRDBUS(98),
	GlitchData    => PPCMPLBWRDBUS98_GlitchData,
	OutSignalName => "PPCMPLBWRDBUS(98)",
	OutTemp       => PPCMPLBWRDBUS_OUT(98),
	Paths         => (0 => (CPMPPCMPLBCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCMPLBWRDBUS(99),
	GlitchData    => PPCMPLBWRDBUS99_GlitchData,
	OutSignalName => "PPCMPLBWRDBUS(99)",
	OutTemp       => PPCMPLBWRDBUS_OUT(99),
	Paths         => (0 => (CPMPPCMPLBCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCMPLBWRDBUS(100),
	GlitchData    => PPCMPLBWRDBUS100_GlitchData,
	OutSignalName => "PPCMPLBWRDBUS(100)",
	OutTemp       => PPCMPLBWRDBUS_OUT(100),
	Paths         => (0 => (CPMPPCMPLBCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCMPLBWRDBUS(101),
	GlitchData    => PPCMPLBWRDBUS101_GlitchData,
	OutSignalName => "PPCMPLBWRDBUS(101)",
	OutTemp       => PPCMPLBWRDBUS_OUT(101),
	Paths         => (0 => (CPMPPCMPLBCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCMPLBWRDBUS(102),
	GlitchData    => PPCMPLBWRDBUS102_GlitchData,
	OutSignalName => "PPCMPLBWRDBUS(102)",
	OutTemp       => PPCMPLBWRDBUS_OUT(102),
	Paths         => (0 => (CPMPPCMPLBCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCMPLBWRDBUS(103),
	GlitchData    => PPCMPLBWRDBUS103_GlitchData,
	OutSignalName => "PPCMPLBWRDBUS(103)",
	OutTemp       => PPCMPLBWRDBUS_OUT(103),
	Paths         => (0 => (CPMPPCMPLBCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCMPLBWRDBUS(104),
	GlitchData    => PPCMPLBWRDBUS104_GlitchData,
	OutSignalName => "PPCMPLBWRDBUS(104)",
	OutTemp       => PPCMPLBWRDBUS_OUT(104),
	Paths         => (0 => (CPMPPCMPLBCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCMPLBWRDBUS(105),
	GlitchData    => PPCMPLBWRDBUS105_GlitchData,
	OutSignalName => "PPCMPLBWRDBUS(105)",
	OutTemp       => PPCMPLBWRDBUS_OUT(105),
	Paths         => (0 => (CPMPPCMPLBCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCMPLBWRDBUS(106),
	GlitchData    => PPCMPLBWRDBUS106_GlitchData,
	OutSignalName => "PPCMPLBWRDBUS(106)",
	OutTemp       => PPCMPLBWRDBUS_OUT(106),
	Paths         => (0 => (CPMPPCMPLBCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCMPLBWRDBUS(107),
	GlitchData    => PPCMPLBWRDBUS107_GlitchData,
	OutSignalName => "PPCMPLBWRDBUS(107)",
	OutTemp       => PPCMPLBWRDBUS_OUT(107),
	Paths         => (0 => (CPMPPCMPLBCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCMPLBWRDBUS(108),
	GlitchData    => PPCMPLBWRDBUS108_GlitchData,
	OutSignalName => "PPCMPLBWRDBUS(108)",
	OutTemp       => PPCMPLBWRDBUS_OUT(108),
	Paths         => (0 => (CPMPPCMPLBCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCMPLBWRDBUS(109),
	GlitchData    => PPCMPLBWRDBUS109_GlitchData,
	OutSignalName => "PPCMPLBWRDBUS(109)",
	OutTemp       => PPCMPLBWRDBUS_OUT(109),
	Paths         => (0 => (CPMPPCMPLBCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCMPLBWRDBUS(110),
	GlitchData    => PPCMPLBWRDBUS110_GlitchData,
	OutSignalName => "PPCMPLBWRDBUS(110)",
	OutTemp       => PPCMPLBWRDBUS_OUT(110),
	Paths         => (0 => (CPMPPCMPLBCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCMPLBWRDBUS(111),
	GlitchData    => PPCMPLBWRDBUS111_GlitchData,
	OutSignalName => "PPCMPLBWRDBUS(111)",
	OutTemp       => PPCMPLBWRDBUS_OUT(111),
	Paths         => (0 => (CPMPPCMPLBCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCMPLBWRDBUS(112),
	GlitchData    => PPCMPLBWRDBUS112_GlitchData,
	OutSignalName => "PPCMPLBWRDBUS(112)",
	OutTemp       => PPCMPLBWRDBUS_OUT(112),
	Paths         => (0 => (CPMPPCMPLBCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCMPLBWRDBUS(113),
	GlitchData    => PPCMPLBWRDBUS113_GlitchData,
	OutSignalName => "PPCMPLBWRDBUS(113)",
	OutTemp       => PPCMPLBWRDBUS_OUT(113),
	Paths         => (0 => (CPMPPCMPLBCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCMPLBWRDBUS(114),
	GlitchData    => PPCMPLBWRDBUS114_GlitchData,
	OutSignalName => "PPCMPLBWRDBUS(114)",
	OutTemp       => PPCMPLBWRDBUS_OUT(114),
	Paths         => (0 => (CPMPPCMPLBCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCMPLBWRDBUS(115),
	GlitchData    => PPCMPLBWRDBUS115_GlitchData,
	OutSignalName => "PPCMPLBWRDBUS(115)",
	OutTemp       => PPCMPLBWRDBUS_OUT(115),
	Paths         => (0 => (CPMPPCMPLBCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCMPLBWRDBUS(116),
	GlitchData    => PPCMPLBWRDBUS116_GlitchData,
	OutSignalName => "PPCMPLBWRDBUS(116)",
	OutTemp       => PPCMPLBWRDBUS_OUT(116),
	Paths         => (0 => (CPMPPCMPLBCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCMPLBWRDBUS(117),
	GlitchData    => PPCMPLBWRDBUS117_GlitchData,
	OutSignalName => "PPCMPLBWRDBUS(117)",
	OutTemp       => PPCMPLBWRDBUS_OUT(117),
	Paths         => (0 => (CPMPPCMPLBCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCMPLBWRDBUS(118),
	GlitchData    => PPCMPLBWRDBUS118_GlitchData,
	OutSignalName => "PPCMPLBWRDBUS(118)",
	OutTemp       => PPCMPLBWRDBUS_OUT(118),
	Paths         => (0 => (CPMPPCMPLBCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCMPLBWRDBUS(119),
	GlitchData    => PPCMPLBWRDBUS119_GlitchData,
	OutSignalName => "PPCMPLBWRDBUS(119)",
	OutTemp       => PPCMPLBWRDBUS_OUT(119),
	Paths         => (0 => (CPMPPCMPLBCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCMPLBWRDBUS(120),
	GlitchData    => PPCMPLBWRDBUS120_GlitchData,
	OutSignalName => "PPCMPLBWRDBUS(120)",
	OutTemp       => PPCMPLBWRDBUS_OUT(120),
	Paths         => (0 => (CPMPPCMPLBCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCMPLBWRDBUS(121),
	GlitchData    => PPCMPLBWRDBUS121_GlitchData,
	OutSignalName => "PPCMPLBWRDBUS(121)",
	OutTemp       => PPCMPLBWRDBUS_OUT(121),
	Paths         => (0 => (CPMPPCMPLBCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCMPLBWRDBUS(122),
	GlitchData    => PPCMPLBWRDBUS122_GlitchData,
	OutSignalName => "PPCMPLBWRDBUS(122)",
	OutTemp       => PPCMPLBWRDBUS_OUT(122),
	Paths         => (0 => (CPMPPCMPLBCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCMPLBWRDBUS(123),
	GlitchData    => PPCMPLBWRDBUS123_GlitchData,
	OutSignalName => "PPCMPLBWRDBUS(123)",
	OutTemp       => PPCMPLBWRDBUS_OUT(123),
	Paths         => (0 => (CPMPPCMPLBCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCMPLBWRDBUS(124),
	GlitchData    => PPCMPLBWRDBUS124_GlitchData,
	OutSignalName => "PPCMPLBWRDBUS(124)",
	OutTemp       => PPCMPLBWRDBUS_OUT(124),
	Paths         => (0 => (CPMPPCMPLBCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCMPLBWRDBUS(125),
	GlitchData    => PPCMPLBWRDBUS125_GlitchData,
	OutSignalName => "PPCMPLBWRDBUS(125)",
	OutTemp       => PPCMPLBWRDBUS_OUT(125),
	Paths         => (0 => (CPMPPCMPLBCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCMPLBWRDBUS(126),
	GlitchData    => PPCMPLBWRDBUS126_GlitchData,
	OutSignalName => "PPCMPLBWRDBUS(126)",
	OutTemp       => PPCMPLBWRDBUS_OUT(126),
	Paths         => (0 => (CPMPPCMPLBCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCMPLBWRDBUS(127),
	GlitchData    => PPCMPLBWRDBUS127_GlitchData,
	OutSignalName => "PPCMPLBWRDBUS(127)",
	OutTemp       => PPCMPLBWRDBUS_OUT(127),
	Paths         => (0 => (CPMPPCMPLBCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS0PLBADDRACK,
	GlitchData    => PPCS0PLBADDRACK_GlitchData,
	OutSignalName => "PPCS0PLBADDRACK",
	OutTemp       => PPCS0PLBADDRACK_OUT,
	Paths         => (0 => (CPMPPCS0PLBCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS0PLBMBUSY(0),
	GlitchData    => PPCS0PLBMBUSY0_GlitchData,
	OutSignalName => "PPCS0PLBMBUSY(0)",
	OutTemp       => PPCS0PLBMBUSY_OUT(0),
	Paths         => (0 => (CPMPPCS0PLBCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS0PLBMBUSY(1),
	GlitchData    => PPCS0PLBMBUSY1_GlitchData,
	OutSignalName => "PPCS0PLBMBUSY(1)",
	OutTemp       => PPCS0PLBMBUSY_OUT(1),
	Paths         => (0 => (CPMPPCS0PLBCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS0PLBMBUSY(2),
	GlitchData    => PPCS0PLBMBUSY2_GlitchData,
	OutSignalName => "PPCS0PLBMBUSY(2)",
	OutTemp       => PPCS0PLBMBUSY_OUT(2),
	Paths         => (0 => (CPMPPCS0PLBCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS0PLBMBUSY(3),
	GlitchData    => PPCS0PLBMBUSY3_GlitchData,
	OutSignalName => "PPCS0PLBMBUSY(3)",
	OutTemp       => PPCS0PLBMBUSY_OUT(3),
	Paths         => (0 => (CPMPPCS0PLBCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS0PLBMIRQ(0),
	GlitchData    => PPCS0PLBMIRQ0_GlitchData,
	OutSignalName => "PPCS0PLBMIRQ(0)",
	OutTemp       => PPCS0PLBMIRQ_OUT(0),
	Paths         => (0 => (CPMPPCS0PLBCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS0PLBMIRQ(1),
	GlitchData    => PPCS0PLBMIRQ1_GlitchData,
	OutSignalName => "PPCS0PLBMIRQ(1)",
	OutTemp       => PPCS0PLBMIRQ_OUT(1),
	Paths         => (0 => (CPMPPCS0PLBCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS0PLBMIRQ(2),
	GlitchData    => PPCS0PLBMIRQ2_GlitchData,
	OutSignalName => "PPCS0PLBMIRQ(2)",
	OutTemp       => PPCS0PLBMIRQ_OUT(2),
	Paths         => (0 => (CPMPPCS0PLBCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS0PLBMIRQ(3),
	GlitchData    => PPCS0PLBMIRQ3_GlitchData,
	OutSignalName => "PPCS0PLBMIRQ(3)",
	OutTemp       => PPCS0PLBMIRQ_OUT(3),
	Paths         => (0 => (CPMPPCS0PLBCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS0PLBMRDERR(0),
	GlitchData    => PPCS0PLBMRDERR0_GlitchData,
	OutSignalName => "PPCS0PLBMRDERR(0)",
	OutTemp       => PPCS0PLBMRDERR_OUT(0),
	Paths         => (0 => (CPMPPCS0PLBCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS0PLBMRDERR(1),
	GlitchData    => PPCS0PLBMRDERR1_GlitchData,
	OutSignalName => "PPCS0PLBMRDERR(1)",
	OutTemp       => PPCS0PLBMRDERR_OUT(1),
	Paths         => (0 => (CPMPPCS0PLBCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS0PLBMRDERR(2),
	GlitchData    => PPCS0PLBMRDERR2_GlitchData,
	OutSignalName => "PPCS0PLBMRDERR(2)",
	OutTemp       => PPCS0PLBMRDERR_OUT(2),
	Paths         => (0 => (CPMPPCS0PLBCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS0PLBMRDERR(3),
	GlitchData    => PPCS0PLBMRDERR3_GlitchData,
	OutSignalName => "PPCS0PLBMRDERR(3)",
	OutTemp       => PPCS0PLBMRDERR_OUT(3),
	Paths         => (0 => (CPMPPCS0PLBCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS0PLBMWRERR(0),
	GlitchData    => PPCS0PLBMWRERR0_GlitchData,
	OutSignalName => "PPCS0PLBMWRERR(0)",
	OutTemp       => PPCS0PLBMWRERR_OUT(0),
	Paths         => (0 => (CPMPPCS0PLBCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS0PLBMWRERR(1),
	GlitchData    => PPCS0PLBMWRERR1_GlitchData,
	OutSignalName => "PPCS0PLBMWRERR(1)",
	OutTemp       => PPCS0PLBMWRERR_OUT(1),
	Paths         => (0 => (CPMPPCS0PLBCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS0PLBMWRERR(2),
	GlitchData    => PPCS0PLBMWRERR2_GlitchData,
	OutSignalName => "PPCS0PLBMWRERR(2)",
	OutTemp       => PPCS0PLBMWRERR_OUT(2),
	Paths         => (0 => (CPMPPCS0PLBCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS0PLBMWRERR(3),
	GlitchData    => PPCS0PLBMWRERR3_GlitchData,
	OutSignalName => "PPCS0PLBMWRERR(3)",
	OutTemp       => PPCS0PLBMWRERR_OUT(3),
	Paths         => (0 => (CPMPPCS0PLBCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS0PLBRDBTERM,
	GlitchData    => PPCS0PLBRDBTERM_GlitchData,
	OutSignalName => "PPCS0PLBRDBTERM",
	OutTemp       => PPCS0PLBRDBTERM_OUT,
	Paths         => (0 => (CPMPPCS0PLBCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS0PLBRDCOMP,
	GlitchData    => PPCS0PLBRDCOMP_GlitchData,
	OutSignalName => "PPCS0PLBRDCOMP",
	OutTemp       => PPCS0PLBRDCOMP_OUT,
	Paths         => (0 => (CPMPPCS0PLBCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS0PLBRDDACK,
	GlitchData    => PPCS0PLBRDDACK_GlitchData,
	OutSignalName => "PPCS0PLBRDDACK",
	OutTemp       => PPCS0PLBRDDACK_OUT,
	Paths         => (0 => (CPMPPCS0PLBCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS0PLBRDDBUS(0),
	GlitchData    => PPCS0PLBRDDBUS0_GlitchData,
	OutSignalName => "PPCS0PLBRDDBUS(0)",
	OutTemp       => PPCS0PLBRDDBUS_OUT(0),
	Paths         => (0 => (CPMPPCS0PLBCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS0PLBRDDBUS(1),
	GlitchData    => PPCS0PLBRDDBUS1_GlitchData,
	OutSignalName => "PPCS0PLBRDDBUS(1)",
	OutTemp       => PPCS0PLBRDDBUS_OUT(1),
	Paths         => (0 => (CPMPPCS0PLBCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS0PLBRDDBUS(2),
	GlitchData    => PPCS0PLBRDDBUS2_GlitchData,
	OutSignalName => "PPCS0PLBRDDBUS(2)",
	OutTemp       => PPCS0PLBRDDBUS_OUT(2),
	Paths         => (0 => (CPMPPCS0PLBCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS0PLBRDDBUS(3),
	GlitchData    => PPCS0PLBRDDBUS3_GlitchData,
	OutSignalName => "PPCS0PLBRDDBUS(3)",
	OutTemp       => PPCS0PLBRDDBUS_OUT(3),
	Paths         => (0 => (CPMPPCS0PLBCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS0PLBRDDBUS(4),
	GlitchData    => PPCS0PLBRDDBUS4_GlitchData,
	OutSignalName => "PPCS0PLBRDDBUS(4)",
	OutTemp       => PPCS0PLBRDDBUS_OUT(4),
	Paths         => (0 => (CPMPPCS0PLBCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS0PLBRDDBUS(5),
	GlitchData    => PPCS0PLBRDDBUS5_GlitchData,
	OutSignalName => "PPCS0PLBRDDBUS(5)",
	OutTemp       => PPCS0PLBRDDBUS_OUT(5),
	Paths         => (0 => (CPMPPCS0PLBCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS0PLBRDDBUS(6),
	GlitchData    => PPCS0PLBRDDBUS6_GlitchData,
	OutSignalName => "PPCS0PLBRDDBUS(6)",
	OutTemp       => PPCS0PLBRDDBUS_OUT(6),
	Paths         => (0 => (CPMPPCS0PLBCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS0PLBRDDBUS(7),
	GlitchData    => PPCS0PLBRDDBUS7_GlitchData,
	OutSignalName => "PPCS0PLBRDDBUS(7)",
	OutTemp       => PPCS0PLBRDDBUS_OUT(7),
	Paths         => (0 => (CPMPPCS0PLBCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS0PLBRDDBUS(8),
	GlitchData    => PPCS0PLBRDDBUS8_GlitchData,
	OutSignalName => "PPCS0PLBRDDBUS(8)",
	OutTemp       => PPCS0PLBRDDBUS_OUT(8),
	Paths         => (0 => (CPMPPCS0PLBCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS0PLBRDDBUS(9),
	GlitchData    => PPCS0PLBRDDBUS9_GlitchData,
	OutSignalName => "PPCS0PLBRDDBUS(9)",
	OutTemp       => PPCS0PLBRDDBUS_OUT(9),
	Paths         => (0 => (CPMPPCS0PLBCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS0PLBRDDBUS(10),
	GlitchData    => PPCS0PLBRDDBUS10_GlitchData,
	OutSignalName => "PPCS0PLBRDDBUS(10)",
	OutTemp       => PPCS0PLBRDDBUS_OUT(10),
	Paths         => (0 => (CPMPPCS0PLBCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS0PLBRDDBUS(11),
	GlitchData    => PPCS0PLBRDDBUS11_GlitchData,
	OutSignalName => "PPCS0PLBRDDBUS(11)",
	OutTemp       => PPCS0PLBRDDBUS_OUT(11),
	Paths         => (0 => (CPMPPCS0PLBCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS0PLBRDDBUS(12),
	GlitchData    => PPCS0PLBRDDBUS12_GlitchData,
	OutSignalName => "PPCS0PLBRDDBUS(12)",
	OutTemp       => PPCS0PLBRDDBUS_OUT(12),
	Paths         => (0 => (CPMPPCS0PLBCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS0PLBRDDBUS(13),
	GlitchData    => PPCS0PLBRDDBUS13_GlitchData,
	OutSignalName => "PPCS0PLBRDDBUS(13)",
	OutTemp       => PPCS0PLBRDDBUS_OUT(13),
	Paths         => (0 => (CPMPPCS0PLBCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS0PLBRDDBUS(14),
	GlitchData    => PPCS0PLBRDDBUS14_GlitchData,
	OutSignalName => "PPCS0PLBRDDBUS(14)",
	OutTemp       => PPCS0PLBRDDBUS_OUT(14),
	Paths         => (0 => (CPMPPCS0PLBCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS0PLBRDDBUS(15),
	GlitchData    => PPCS0PLBRDDBUS15_GlitchData,
	OutSignalName => "PPCS0PLBRDDBUS(15)",
	OutTemp       => PPCS0PLBRDDBUS_OUT(15),
	Paths         => (0 => (CPMPPCS0PLBCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS0PLBRDDBUS(16),
	GlitchData    => PPCS0PLBRDDBUS16_GlitchData,
	OutSignalName => "PPCS0PLBRDDBUS(16)",
	OutTemp       => PPCS0PLBRDDBUS_OUT(16),
	Paths         => (0 => (CPMPPCS0PLBCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS0PLBRDDBUS(17),
	GlitchData    => PPCS0PLBRDDBUS17_GlitchData,
	OutSignalName => "PPCS0PLBRDDBUS(17)",
	OutTemp       => PPCS0PLBRDDBUS_OUT(17),
	Paths         => (0 => (CPMPPCS0PLBCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS0PLBRDDBUS(18),
	GlitchData    => PPCS0PLBRDDBUS18_GlitchData,
	OutSignalName => "PPCS0PLBRDDBUS(18)",
	OutTemp       => PPCS0PLBRDDBUS_OUT(18),
	Paths         => (0 => (CPMPPCS0PLBCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS0PLBRDDBUS(19),
	GlitchData    => PPCS0PLBRDDBUS19_GlitchData,
	OutSignalName => "PPCS0PLBRDDBUS(19)",
	OutTemp       => PPCS0PLBRDDBUS_OUT(19),
	Paths         => (0 => (CPMPPCS0PLBCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS0PLBRDDBUS(20),
	GlitchData    => PPCS0PLBRDDBUS20_GlitchData,
	OutSignalName => "PPCS0PLBRDDBUS(20)",
	OutTemp       => PPCS0PLBRDDBUS_OUT(20),
	Paths         => (0 => (CPMPPCS0PLBCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS0PLBRDDBUS(21),
	GlitchData    => PPCS0PLBRDDBUS21_GlitchData,
	OutSignalName => "PPCS0PLBRDDBUS(21)",
	OutTemp       => PPCS0PLBRDDBUS_OUT(21),
	Paths         => (0 => (CPMPPCS0PLBCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS0PLBRDDBUS(22),
	GlitchData    => PPCS0PLBRDDBUS22_GlitchData,
	OutSignalName => "PPCS0PLBRDDBUS(22)",
	OutTemp       => PPCS0PLBRDDBUS_OUT(22),
	Paths         => (0 => (CPMPPCS0PLBCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS0PLBRDDBUS(23),
	GlitchData    => PPCS0PLBRDDBUS23_GlitchData,
	OutSignalName => "PPCS0PLBRDDBUS(23)",
	OutTemp       => PPCS0PLBRDDBUS_OUT(23),
	Paths         => (0 => (CPMPPCS0PLBCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS0PLBRDDBUS(24),
	GlitchData    => PPCS0PLBRDDBUS24_GlitchData,
	OutSignalName => "PPCS0PLBRDDBUS(24)",
	OutTemp       => PPCS0PLBRDDBUS_OUT(24),
	Paths         => (0 => (CPMPPCS0PLBCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS0PLBRDDBUS(25),
	GlitchData    => PPCS0PLBRDDBUS25_GlitchData,
	OutSignalName => "PPCS0PLBRDDBUS(25)",
	OutTemp       => PPCS0PLBRDDBUS_OUT(25),
	Paths         => (0 => (CPMPPCS0PLBCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS0PLBRDDBUS(26),
	GlitchData    => PPCS0PLBRDDBUS26_GlitchData,
	OutSignalName => "PPCS0PLBRDDBUS(26)",
	OutTemp       => PPCS0PLBRDDBUS_OUT(26),
	Paths         => (0 => (CPMPPCS0PLBCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS0PLBRDDBUS(27),
	GlitchData    => PPCS0PLBRDDBUS27_GlitchData,
	OutSignalName => "PPCS0PLBRDDBUS(27)",
	OutTemp       => PPCS0PLBRDDBUS_OUT(27),
	Paths         => (0 => (CPMPPCS0PLBCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS0PLBRDDBUS(28),
	GlitchData    => PPCS0PLBRDDBUS28_GlitchData,
	OutSignalName => "PPCS0PLBRDDBUS(28)",
	OutTemp       => PPCS0PLBRDDBUS_OUT(28),
	Paths         => (0 => (CPMPPCS0PLBCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS0PLBRDDBUS(29),
	GlitchData    => PPCS0PLBRDDBUS29_GlitchData,
	OutSignalName => "PPCS0PLBRDDBUS(29)",
	OutTemp       => PPCS0PLBRDDBUS_OUT(29),
	Paths         => (0 => (CPMPPCS0PLBCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS0PLBRDDBUS(30),
	GlitchData    => PPCS0PLBRDDBUS30_GlitchData,
	OutSignalName => "PPCS0PLBRDDBUS(30)",
	OutTemp       => PPCS0PLBRDDBUS_OUT(30),
	Paths         => (0 => (CPMPPCS0PLBCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS0PLBRDDBUS(31),
	GlitchData    => PPCS0PLBRDDBUS31_GlitchData,
	OutSignalName => "PPCS0PLBRDDBUS(31)",
	OutTemp       => PPCS0PLBRDDBUS_OUT(31),
	Paths         => (0 => (CPMPPCS0PLBCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS0PLBRDDBUS(32),
	GlitchData    => PPCS0PLBRDDBUS32_GlitchData,
	OutSignalName => "PPCS0PLBRDDBUS(32)",
	OutTemp       => PPCS0PLBRDDBUS_OUT(32),
	Paths         => (0 => (CPMPPCS0PLBCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS0PLBRDDBUS(33),
	GlitchData    => PPCS0PLBRDDBUS33_GlitchData,
	OutSignalName => "PPCS0PLBRDDBUS(33)",
	OutTemp       => PPCS0PLBRDDBUS_OUT(33),
	Paths         => (0 => (CPMPPCS0PLBCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS0PLBRDDBUS(34),
	GlitchData    => PPCS0PLBRDDBUS34_GlitchData,
	OutSignalName => "PPCS0PLBRDDBUS(34)",
	OutTemp       => PPCS0PLBRDDBUS_OUT(34),
	Paths         => (0 => (CPMPPCS0PLBCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS0PLBRDDBUS(35),
	GlitchData    => PPCS0PLBRDDBUS35_GlitchData,
	OutSignalName => "PPCS0PLBRDDBUS(35)",
	OutTemp       => PPCS0PLBRDDBUS_OUT(35),
	Paths         => (0 => (CPMPPCS0PLBCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS0PLBRDDBUS(36),
	GlitchData    => PPCS0PLBRDDBUS36_GlitchData,
	OutSignalName => "PPCS0PLBRDDBUS(36)",
	OutTemp       => PPCS0PLBRDDBUS_OUT(36),
	Paths         => (0 => (CPMPPCS0PLBCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS0PLBRDDBUS(37),
	GlitchData    => PPCS0PLBRDDBUS37_GlitchData,
	OutSignalName => "PPCS0PLBRDDBUS(37)",
	OutTemp       => PPCS0PLBRDDBUS_OUT(37),
	Paths         => (0 => (CPMPPCS0PLBCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS0PLBRDDBUS(38),
	GlitchData    => PPCS0PLBRDDBUS38_GlitchData,
	OutSignalName => "PPCS0PLBRDDBUS(38)",
	OutTemp       => PPCS0PLBRDDBUS_OUT(38),
	Paths         => (0 => (CPMPPCS0PLBCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS0PLBRDDBUS(39),
	GlitchData    => PPCS0PLBRDDBUS39_GlitchData,
	OutSignalName => "PPCS0PLBRDDBUS(39)",
	OutTemp       => PPCS0PLBRDDBUS_OUT(39),
	Paths         => (0 => (CPMPPCS0PLBCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS0PLBRDDBUS(40),
	GlitchData    => PPCS0PLBRDDBUS40_GlitchData,
	OutSignalName => "PPCS0PLBRDDBUS(40)",
	OutTemp       => PPCS0PLBRDDBUS_OUT(40),
	Paths         => (0 => (CPMPPCS0PLBCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS0PLBRDDBUS(41),
	GlitchData    => PPCS0PLBRDDBUS41_GlitchData,
	OutSignalName => "PPCS0PLBRDDBUS(41)",
	OutTemp       => PPCS0PLBRDDBUS_OUT(41),
	Paths         => (0 => (CPMPPCS0PLBCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS0PLBRDDBUS(42),
	GlitchData    => PPCS0PLBRDDBUS42_GlitchData,
	OutSignalName => "PPCS0PLBRDDBUS(42)",
	OutTemp       => PPCS0PLBRDDBUS_OUT(42),
	Paths         => (0 => (CPMPPCS0PLBCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS0PLBRDDBUS(43),
	GlitchData    => PPCS0PLBRDDBUS43_GlitchData,
	OutSignalName => "PPCS0PLBRDDBUS(43)",
	OutTemp       => PPCS0PLBRDDBUS_OUT(43),
	Paths         => (0 => (CPMPPCS0PLBCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS0PLBRDDBUS(44),
	GlitchData    => PPCS0PLBRDDBUS44_GlitchData,
	OutSignalName => "PPCS0PLBRDDBUS(44)",
	OutTemp       => PPCS0PLBRDDBUS_OUT(44),
	Paths         => (0 => (CPMPPCS0PLBCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS0PLBRDDBUS(45),
	GlitchData    => PPCS0PLBRDDBUS45_GlitchData,
	OutSignalName => "PPCS0PLBRDDBUS(45)",
	OutTemp       => PPCS0PLBRDDBUS_OUT(45),
	Paths         => (0 => (CPMPPCS0PLBCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS0PLBRDDBUS(46),
	GlitchData    => PPCS0PLBRDDBUS46_GlitchData,
	OutSignalName => "PPCS0PLBRDDBUS(46)",
	OutTemp       => PPCS0PLBRDDBUS_OUT(46),
	Paths         => (0 => (CPMPPCS0PLBCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS0PLBRDDBUS(47),
	GlitchData    => PPCS0PLBRDDBUS47_GlitchData,
	OutSignalName => "PPCS0PLBRDDBUS(47)",
	OutTemp       => PPCS0PLBRDDBUS_OUT(47),
	Paths         => (0 => (CPMPPCS0PLBCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS0PLBRDDBUS(48),
	GlitchData    => PPCS0PLBRDDBUS48_GlitchData,
	OutSignalName => "PPCS0PLBRDDBUS(48)",
	OutTemp       => PPCS0PLBRDDBUS_OUT(48),
	Paths         => (0 => (CPMPPCS0PLBCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS0PLBRDDBUS(49),
	GlitchData    => PPCS0PLBRDDBUS49_GlitchData,
	OutSignalName => "PPCS0PLBRDDBUS(49)",
	OutTemp       => PPCS0PLBRDDBUS_OUT(49),
	Paths         => (0 => (CPMPPCS0PLBCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS0PLBRDDBUS(50),
	GlitchData    => PPCS0PLBRDDBUS50_GlitchData,
	OutSignalName => "PPCS0PLBRDDBUS(50)",
	OutTemp       => PPCS0PLBRDDBUS_OUT(50),
	Paths         => (0 => (CPMPPCS0PLBCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS0PLBRDDBUS(51),
	GlitchData    => PPCS0PLBRDDBUS51_GlitchData,
	OutSignalName => "PPCS0PLBRDDBUS(51)",
	OutTemp       => PPCS0PLBRDDBUS_OUT(51),
	Paths         => (0 => (CPMPPCS0PLBCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS0PLBRDDBUS(52),
	GlitchData    => PPCS0PLBRDDBUS52_GlitchData,
	OutSignalName => "PPCS0PLBRDDBUS(52)",
	OutTemp       => PPCS0PLBRDDBUS_OUT(52),
	Paths         => (0 => (CPMPPCS0PLBCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS0PLBRDDBUS(53),
	GlitchData    => PPCS0PLBRDDBUS53_GlitchData,
	OutSignalName => "PPCS0PLBRDDBUS(53)",
	OutTemp       => PPCS0PLBRDDBUS_OUT(53),
	Paths         => (0 => (CPMPPCS0PLBCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS0PLBRDDBUS(54),
	GlitchData    => PPCS0PLBRDDBUS54_GlitchData,
	OutSignalName => "PPCS0PLBRDDBUS(54)",
	OutTemp       => PPCS0PLBRDDBUS_OUT(54),
	Paths         => (0 => (CPMPPCS0PLBCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS0PLBRDDBUS(55),
	GlitchData    => PPCS0PLBRDDBUS55_GlitchData,
	OutSignalName => "PPCS0PLBRDDBUS(55)",
	OutTemp       => PPCS0PLBRDDBUS_OUT(55),
	Paths         => (0 => (CPMPPCS0PLBCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS0PLBRDDBUS(56),
	GlitchData    => PPCS0PLBRDDBUS56_GlitchData,
	OutSignalName => "PPCS0PLBRDDBUS(56)",
	OutTemp       => PPCS0PLBRDDBUS_OUT(56),
	Paths         => (0 => (CPMPPCS0PLBCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS0PLBRDDBUS(57),
	GlitchData    => PPCS0PLBRDDBUS57_GlitchData,
	OutSignalName => "PPCS0PLBRDDBUS(57)",
	OutTemp       => PPCS0PLBRDDBUS_OUT(57),
	Paths         => (0 => (CPMPPCS0PLBCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS0PLBRDDBUS(58),
	GlitchData    => PPCS0PLBRDDBUS58_GlitchData,
	OutSignalName => "PPCS0PLBRDDBUS(58)",
	OutTemp       => PPCS0PLBRDDBUS_OUT(58),
	Paths         => (0 => (CPMPPCS0PLBCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS0PLBRDDBUS(59),
	GlitchData    => PPCS0PLBRDDBUS59_GlitchData,
	OutSignalName => "PPCS0PLBRDDBUS(59)",
	OutTemp       => PPCS0PLBRDDBUS_OUT(59),
	Paths         => (0 => (CPMPPCS0PLBCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS0PLBRDDBUS(60),
	GlitchData    => PPCS0PLBRDDBUS60_GlitchData,
	OutSignalName => "PPCS0PLBRDDBUS(60)",
	OutTemp       => PPCS0PLBRDDBUS_OUT(60),
	Paths         => (0 => (CPMPPCS0PLBCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS0PLBRDDBUS(61),
	GlitchData    => PPCS0PLBRDDBUS61_GlitchData,
	OutSignalName => "PPCS0PLBRDDBUS(61)",
	OutTemp       => PPCS0PLBRDDBUS_OUT(61),
	Paths         => (0 => (CPMPPCS0PLBCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS0PLBRDDBUS(62),
	GlitchData    => PPCS0PLBRDDBUS62_GlitchData,
	OutSignalName => "PPCS0PLBRDDBUS(62)",
	OutTemp       => PPCS0PLBRDDBUS_OUT(62),
	Paths         => (0 => (CPMPPCS0PLBCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS0PLBRDDBUS(63),
	GlitchData    => PPCS0PLBRDDBUS63_GlitchData,
	OutSignalName => "PPCS0PLBRDDBUS(63)",
	OutTemp       => PPCS0PLBRDDBUS_OUT(63),
	Paths         => (0 => (CPMPPCS0PLBCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS0PLBRDDBUS(64),
	GlitchData    => PPCS0PLBRDDBUS64_GlitchData,
	OutSignalName => "PPCS0PLBRDDBUS(64)",
	OutTemp       => PPCS0PLBRDDBUS_OUT(64),
	Paths         => (0 => (CPMPPCS0PLBCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS0PLBRDDBUS(65),
	GlitchData    => PPCS0PLBRDDBUS65_GlitchData,
	OutSignalName => "PPCS0PLBRDDBUS(65)",
	OutTemp       => PPCS0PLBRDDBUS_OUT(65),
	Paths         => (0 => (CPMPPCS0PLBCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS0PLBRDDBUS(66),
	GlitchData    => PPCS0PLBRDDBUS66_GlitchData,
	OutSignalName => "PPCS0PLBRDDBUS(66)",
	OutTemp       => PPCS0PLBRDDBUS_OUT(66),
	Paths         => (0 => (CPMPPCS0PLBCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS0PLBRDDBUS(67),
	GlitchData    => PPCS0PLBRDDBUS67_GlitchData,
	OutSignalName => "PPCS0PLBRDDBUS(67)",
	OutTemp       => PPCS0PLBRDDBUS_OUT(67),
	Paths         => (0 => (CPMPPCS0PLBCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS0PLBRDDBUS(68),
	GlitchData    => PPCS0PLBRDDBUS68_GlitchData,
	OutSignalName => "PPCS0PLBRDDBUS(68)",
	OutTemp       => PPCS0PLBRDDBUS_OUT(68),
	Paths         => (0 => (CPMPPCS0PLBCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS0PLBRDDBUS(69),
	GlitchData    => PPCS0PLBRDDBUS69_GlitchData,
	OutSignalName => "PPCS0PLBRDDBUS(69)",
	OutTemp       => PPCS0PLBRDDBUS_OUT(69),
	Paths         => (0 => (CPMPPCS0PLBCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS0PLBRDDBUS(70),
	GlitchData    => PPCS0PLBRDDBUS70_GlitchData,
	OutSignalName => "PPCS0PLBRDDBUS(70)",
	OutTemp       => PPCS0PLBRDDBUS_OUT(70),
	Paths         => (0 => (CPMPPCS0PLBCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS0PLBRDDBUS(71),
	GlitchData    => PPCS0PLBRDDBUS71_GlitchData,
	OutSignalName => "PPCS0PLBRDDBUS(71)",
	OutTemp       => PPCS0PLBRDDBUS_OUT(71),
	Paths         => (0 => (CPMPPCS0PLBCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS0PLBRDDBUS(72),
	GlitchData    => PPCS0PLBRDDBUS72_GlitchData,
	OutSignalName => "PPCS0PLBRDDBUS(72)",
	OutTemp       => PPCS0PLBRDDBUS_OUT(72),
	Paths         => (0 => (CPMPPCS0PLBCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS0PLBRDDBUS(73),
	GlitchData    => PPCS0PLBRDDBUS73_GlitchData,
	OutSignalName => "PPCS0PLBRDDBUS(73)",
	OutTemp       => PPCS0PLBRDDBUS_OUT(73),
	Paths         => (0 => (CPMPPCS0PLBCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS0PLBRDDBUS(74),
	GlitchData    => PPCS0PLBRDDBUS74_GlitchData,
	OutSignalName => "PPCS0PLBRDDBUS(74)",
	OutTemp       => PPCS0PLBRDDBUS_OUT(74),
	Paths         => (0 => (CPMPPCS0PLBCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS0PLBRDDBUS(75),
	GlitchData    => PPCS0PLBRDDBUS75_GlitchData,
	OutSignalName => "PPCS0PLBRDDBUS(75)",
	OutTemp       => PPCS0PLBRDDBUS_OUT(75),
	Paths         => (0 => (CPMPPCS0PLBCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS0PLBRDDBUS(76),
	GlitchData    => PPCS0PLBRDDBUS76_GlitchData,
	OutSignalName => "PPCS0PLBRDDBUS(76)",
	OutTemp       => PPCS0PLBRDDBUS_OUT(76),
	Paths         => (0 => (CPMPPCS0PLBCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS0PLBRDDBUS(77),
	GlitchData    => PPCS0PLBRDDBUS77_GlitchData,
	OutSignalName => "PPCS0PLBRDDBUS(77)",
	OutTemp       => PPCS0PLBRDDBUS_OUT(77),
	Paths         => (0 => (CPMPPCS0PLBCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS0PLBRDDBUS(78),
	GlitchData    => PPCS0PLBRDDBUS78_GlitchData,
	OutSignalName => "PPCS0PLBRDDBUS(78)",
	OutTemp       => PPCS0PLBRDDBUS_OUT(78),
	Paths         => (0 => (CPMPPCS0PLBCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS0PLBRDDBUS(79),
	GlitchData    => PPCS0PLBRDDBUS79_GlitchData,
	OutSignalName => "PPCS0PLBRDDBUS(79)",
	OutTemp       => PPCS0PLBRDDBUS_OUT(79),
	Paths         => (0 => (CPMPPCS0PLBCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS0PLBRDDBUS(80),
	GlitchData    => PPCS0PLBRDDBUS80_GlitchData,
	OutSignalName => "PPCS0PLBRDDBUS(80)",
	OutTemp       => PPCS0PLBRDDBUS_OUT(80),
	Paths         => (0 => (CPMPPCS0PLBCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS0PLBRDDBUS(81),
	GlitchData    => PPCS0PLBRDDBUS81_GlitchData,
	OutSignalName => "PPCS0PLBRDDBUS(81)",
	OutTemp       => PPCS0PLBRDDBUS_OUT(81),
	Paths         => (0 => (CPMPPCS0PLBCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS0PLBRDDBUS(82),
	GlitchData    => PPCS0PLBRDDBUS82_GlitchData,
	OutSignalName => "PPCS0PLBRDDBUS(82)",
	OutTemp       => PPCS0PLBRDDBUS_OUT(82),
	Paths         => (0 => (CPMPPCS0PLBCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS0PLBRDDBUS(83),
	GlitchData    => PPCS0PLBRDDBUS83_GlitchData,
	OutSignalName => "PPCS0PLBRDDBUS(83)",
	OutTemp       => PPCS0PLBRDDBUS_OUT(83),
	Paths         => (0 => (CPMPPCS0PLBCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS0PLBRDDBUS(84),
	GlitchData    => PPCS0PLBRDDBUS84_GlitchData,
	OutSignalName => "PPCS0PLBRDDBUS(84)",
	OutTemp       => PPCS0PLBRDDBUS_OUT(84),
	Paths         => (0 => (CPMPPCS0PLBCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS0PLBRDDBUS(85),
	GlitchData    => PPCS0PLBRDDBUS85_GlitchData,
	OutSignalName => "PPCS0PLBRDDBUS(85)",
	OutTemp       => PPCS0PLBRDDBUS_OUT(85),
	Paths         => (0 => (CPMPPCS0PLBCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS0PLBRDDBUS(86),
	GlitchData    => PPCS0PLBRDDBUS86_GlitchData,
	OutSignalName => "PPCS0PLBRDDBUS(86)",
	OutTemp       => PPCS0PLBRDDBUS_OUT(86),
	Paths         => (0 => (CPMPPCS0PLBCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS0PLBRDDBUS(87),
	GlitchData    => PPCS0PLBRDDBUS87_GlitchData,
	OutSignalName => "PPCS0PLBRDDBUS(87)",
	OutTemp       => PPCS0PLBRDDBUS_OUT(87),
	Paths         => (0 => (CPMPPCS0PLBCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS0PLBRDDBUS(88),
	GlitchData    => PPCS0PLBRDDBUS88_GlitchData,
	OutSignalName => "PPCS0PLBRDDBUS(88)",
	OutTemp       => PPCS0PLBRDDBUS_OUT(88),
	Paths         => (0 => (CPMPPCS0PLBCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS0PLBRDDBUS(89),
	GlitchData    => PPCS0PLBRDDBUS89_GlitchData,
	OutSignalName => "PPCS0PLBRDDBUS(89)",
	OutTemp       => PPCS0PLBRDDBUS_OUT(89),
	Paths         => (0 => (CPMPPCS0PLBCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS0PLBRDDBUS(90),
	GlitchData    => PPCS0PLBRDDBUS90_GlitchData,
	OutSignalName => "PPCS0PLBRDDBUS(90)",
	OutTemp       => PPCS0PLBRDDBUS_OUT(90),
	Paths         => (0 => (CPMPPCS0PLBCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS0PLBRDDBUS(91),
	GlitchData    => PPCS0PLBRDDBUS91_GlitchData,
	OutSignalName => "PPCS0PLBRDDBUS(91)",
	OutTemp       => PPCS0PLBRDDBUS_OUT(91),
	Paths         => (0 => (CPMPPCS0PLBCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS0PLBRDDBUS(92),
	GlitchData    => PPCS0PLBRDDBUS92_GlitchData,
	OutSignalName => "PPCS0PLBRDDBUS(92)",
	OutTemp       => PPCS0PLBRDDBUS_OUT(92),
	Paths         => (0 => (CPMPPCS0PLBCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS0PLBRDDBUS(93),
	GlitchData    => PPCS0PLBRDDBUS93_GlitchData,
	OutSignalName => "PPCS0PLBRDDBUS(93)",
	OutTemp       => PPCS0PLBRDDBUS_OUT(93),
	Paths         => (0 => (CPMPPCS0PLBCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS0PLBRDDBUS(94),
	GlitchData    => PPCS0PLBRDDBUS94_GlitchData,
	OutSignalName => "PPCS0PLBRDDBUS(94)",
	OutTemp       => PPCS0PLBRDDBUS_OUT(94),
	Paths         => (0 => (CPMPPCS0PLBCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS0PLBRDDBUS(95),
	GlitchData    => PPCS0PLBRDDBUS95_GlitchData,
	OutSignalName => "PPCS0PLBRDDBUS(95)",
	OutTemp       => PPCS0PLBRDDBUS_OUT(95),
	Paths         => (0 => (CPMPPCS0PLBCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS0PLBRDDBUS(96),
	GlitchData    => PPCS0PLBRDDBUS96_GlitchData,
	OutSignalName => "PPCS0PLBRDDBUS(96)",
	OutTemp       => PPCS0PLBRDDBUS_OUT(96),
	Paths         => (0 => (CPMPPCS0PLBCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS0PLBRDDBUS(97),
	GlitchData    => PPCS0PLBRDDBUS97_GlitchData,
	OutSignalName => "PPCS0PLBRDDBUS(97)",
	OutTemp       => PPCS0PLBRDDBUS_OUT(97),
	Paths         => (0 => (CPMPPCS0PLBCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS0PLBRDDBUS(98),
	GlitchData    => PPCS0PLBRDDBUS98_GlitchData,
	OutSignalName => "PPCS0PLBRDDBUS(98)",
	OutTemp       => PPCS0PLBRDDBUS_OUT(98),
	Paths         => (0 => (CPMPPCS0PLBCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS0PLBRDDBUS(99),
	GlitchData    => PPCS0PLBRDDBUS99_GlitchData,
	OutSignalName => "PPCS0PLBRDDBUS(99)",
	OutTemp       => PPCS0PLBRDDBUS_OUT(99),
	Paths         => (0 => (CPMPPCS0PLBCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS0PLBRDDBUS(100),
	GlitchData    => PPCS0PLBRDDBUS100_GlitchData,
	OutSignalName => "PPCS0PLBRDDBUS(100)",
	OutTemp       => PPCS0PLBRDDBUS_OUT(100),
	Paths         => (0 => (CPMPPCS0PLBCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS0PLBRDDBUS(101),
	GlitchData    => PPCS0PLBRDDBUS101_GlitchData,
	OutSignalName => "PPCS0PLBRDDBUS(101)",
	OutTemp       => PPCS0PLBRDDBUS_OUT(101),
	Paths         => (0 => (CPMPPCS0PLBCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS0PLBRDDBUS(102),
	GlitchData    => PPCS0PLBRDDBUS102_GlitchData,
	OutSignalName => "PPCS0PLBRDDBUS(102)",
	OutTemp       => PPCS0PLBRDDBUS_OUT(102),
	Paths         => (0 => (CPMPPCS0PLBCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS0PLBRDDBUS(103),
	GlitchData    => PPCS0PLBRDDBUS103_GlitchData,
	OutSignalName => "PPCS0PLBRDDBUS(103)",
	OutTemp       => PPCS0PLBRDDBUS_OUT(103),
	Paths         => (0 => (CPMPPCS0PLBCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS0PLBRDDBUS(104),
	GlitchData    => PPCS0PLBRDDBUS104_GlitchData,
	OutSignalName => "PPCS0PLBRDDBUS(104)",
	OutTemp       => PPCS0PLBRDDBUS_OUT(104),
	Paths         => (0 => (CPMPPCS0PLBCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS0PLBRDDBUS(105),
	GlitchData    => PPCS0PLBRDDBUS105_GlitchData,
	OutSignalName => "PPCS0PLBRDDBUS(105)",
	OutTemp       => PPCS0PLBRDDBUS_OUT(105),
	Paths         => (0 => (CPMPPCS0PLBCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS0PLBRDDBUS(106),
	GlitchData    => PPCS0PLBRDDBUS106_GlitchData,
	OutSignalName => "PPCS0PLBRDDBUS(106)",
	OutTemp       => PPCS0PLBRDDBUS_OUT(106),
	Paths         => (0 => (CPMPPCS0PLBCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS0PLBRDDBUS(107),
	GlitchData    => PPCS0PLBRDDBUS107_GlitchData,
	OutSignalName => "PPCS0PLBRDDBUS(107)",
	OutTemp       => PPCS0PLBRDDBUS_OUT(107),
	Paths         => (0 => (CPMPPCS0PLBCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS0PLBRDDBUS(108),
	GlitchData    => PPCS0PLBRDDBUS108_GlitchData,
	OutSignalName => "PPCS0PLBRDDBUS(108)",
	OutTemp       => PPCS0PLBRDDBUS_OUT(108),
	Paths         => (0 => (CPMPPCS0PLBCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS0PLBRDDBUS(109),
	GlitchData    => PPCS0PLBRDDBUS109_GlitchData,
	OutSignalName => "PPCS0PLBRDDBUS(109)",
	OutTemp       => PPCS0PLBRDDBUS_OUT(109),
	Paths         => (0 => (CPMPPCS0PLBCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS0PLBRDDBUS(110),
	GlitchData    => PPCS0PLBRDDBUS110_GlitchData,
	OutSignalName => "PPCS0PLBRDDBUS(110)",
	OutTemp       => PPCS0PLBRDDBUS_OUT(110),
	Paths         => (0 => (CPMPPCS0PLBCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS0PLBRDDBUS(111),
	GlitchData    => PPCS0PLBRDDBUS111_GlitchData,
	OutSignalName => "PPCS0PLBRDDBUS(111)",
	OutTemp       => PPCS0PLBRDDBUS_OUT(111),
	Paths         => (0 => (CPMPPCS0PLBCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS0PLBRDDBUS(112),
	GlitchData    => PPCS0PLBRDDBUS112_GlitchData,
	OutSignalName => "PPCS0PLBRDDBUS(112)",
	OutTemp       => PPCS0PLBRDDBUS_OUT(112),
	Paths         => (0 => (CPMPPCS0PLBCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS0PLBRDDBUS(113),
	GlitchData    => PPCS0PLBRDDBUS113_GlitchData,
	OutSignalName => "PPCS0PLBRDDBUS(113)",
	OutTemp       => PPCS0PLBRDDBUS_OUT(113),
	Paths         => (0 => (CPMPPCS0PLBCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS0PLBRDDBUS(114),
	GlitchData    => PPCS0PLBRDDBUS114_GlitchData,
	OutSignalName => "PPCS0PLBRDDBUS(114)",
	OutTemp       => PPCS0PLBRDDBUS_OUT(114),
	Paths         => (0 => (CPMPPCS0PLBCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS0PLBRDDBUS(115),
	GlitchData    => PPCS0PLBRDDBUS115_GlitchData,
	OutSignalName => "PPCS0PLBRDDBUS(115)",
	OutTemp       => PPCS0PLBRDDBUS_OUT(115),
	Paths         => (0 => (CPMPPCS0PLBCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS0PLBRDDBUS(116),
	GlitchData    => PPCS0PLBRDDBUS116_GlitchData,
	OutSignalName => "PPCS0PLBRDDBUS(116)",
	OutTemp       => PPCS0PLBRDDBUS_OUT(116),
	Paths         => (0 => (CPMPPCS0PLBCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS0PLBRDDBUS(117),
	GlitchData    => PPCS0PLBRDDBUS117_GlitchData,
	OutSignalName => "PPCS0PLBRDDBUS(117)",
	OutTemp       => PPCS0PLBRDDBUS_OUT(117),
	Paths         => (0 => (CPMPPCS0PLBCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS0PLBRDDBUS(118),
	GlitchData    => PPCS0PLBRDDBUS118_GlitchData,
	OutSignalName => "PPCS0PLBRDDBUS(118)",
	OutTemp       => PPCS0PLBRDDBUS_OUT(118),
	Paths         => (0 => (CPMPPCS0PLBCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS0PLBRDDBUS(119),
	GlitchData    => PPCS0PLBRDDBUS119_GlitchData,
	OutSignalName => "PPCS0PLBRDDBUS(119)",
	OutTemp       => PPCS0PLBRDDBUS_OUT(119),
	Paths         => (0 => (CPMPPCS0PLBCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS0PLBRDDBUS(120),
	GlitchData    => PPCS0PLBRDDBUS120_GlitchData,
	OutSignalName => "PPCS0PLBRDDBUS(120)",
	OutTemp       => PPCS0PLBRDDBUS_OUT(120),
	Paths         => (0 => (CPMPPCS0PLBCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS0PLBRDDBUS(121),
	GlitchData    => PPCS0PLBRDDBUS121_GlitchData,
	OutSignalName => "PPCS0PLBRDDBUS(121)",
	OutTemp       => PPCS0PLBRDDBUS_OUT(121),
	Paths         => (0 => (CPMPPCS0PLBCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS0PLBRDDBUS(122),
	GlitchData    => PPCS0PLBRDDBUS122_GlitchData,
	OutSignalName => "PPCS0PLBRDDBUS(122)",
	OutTemp       => PPCS0PLBRDDBUS_OUT(122),
	Paths         => (0 => (CPMPPCS0PLBCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS0PLBRDDBUS(123),
	GlitchData    => PPCS0PLBRDDBUS123_GlitchData,
	OutSignalName => "PPCS0PLBRDDBUS(123)",
	OutTemp       => PPCS0PLBRDDBUS_OUT(123),
	Paths         => (0 => (CPMPPCS0PLBCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS0PLBRDDBUS(124),
	GlitchData    => PPCS0PLBRDDBUS124_GlitchData,
	OutSignalName => "PPCS0PLBRDDBUS(124)",
	OutTemp       => PPCS0PLBRDDBUS_OUT(124),
	Paths         => (0 => (CPMPPCS0PLBCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS0PLBRDDBUS(125),
	GlitchData    => PPCS0PLBRDDBUS125_GlitchData,
	OutSignalName => "PPCS0PLBRDDBUS(125)",
	OutTemp       => PPCS0PLBRDDBUS_OUT(125),
	Paths         => (0 => (CPMPPCS0PLBCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS0PLBRDDBUS(126),
	GlitchData    => PPCS0PLBRDDBUS126_GlitchData,
	OutSignalName => "PPCS0PLBRDDBUS(126)",
	OutTemp       => PPCS0PLBRDDBUS_OUT(126),
	Paths         => (0 => (CPMPPCS0PLBCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS0PLBRDDBUS(127),
	GlitchData    => PPCS0PLBRDDBUS127_GlitchData,
	OutSignalName => "PPCS0PLBRDDBUS(127)",
	OutTemp       => PPCS0PLBRDDBUS_OUT(127),
	Paths         => (0 => (CPMPPCS0PLBCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS0PLBRDWDADDR(0),
	GlitchData    => PPCS0PLBRDWDADDR0_GlitchData,
	OutSignalName => "PPCS0PLBRDWDADDR(0)",
	OutTemp       => PPCS0PLBRDWDADDR_OUT(0),
	Paths         => (0 => (CPMPPCS0PLBCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS0PLBRDWDADDR(1),
	GlitchData    => PPCS0PLBRDWDADDR1_GlitchData,
	OutSignalName => "PPCS0PLBRDWDADDR(1)",
	OutTemp       => PPCS0PLBRDWDADDR_OUT(1),
	Paths         => (0 => (CPMPPCS0PLBCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS0PLBRDWDADDR(2),
	GlitchData    => PPCS0PLBRDWDADDR2_GlitchData,
	OutSignalName => "PPCS0PLBRDWDADDR(2)",
	OutTemp       => PPCS0PLBRDWDADDR_OUT(2),
	Paths         => (0 => (CPMPPCS0PLBCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS0PLBRDWDADDR(3),
	GlitchData    => PPCS0PLBRDWDADDR3_GlitchData,
	OutSignalName => "PPCS0PLBRDWDADDR(3)",
	OutTemp       => PPCS0PLBRDWDADDR_OUT(3),
	Paths         => (0 => (CPMPPCS0PLBCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS0PLBREARBITRATE,
	GlitchData    => PPCS0PLBREARBITRATE_GlitchData,
	OutSignalName => "PPCS0PLBREARBITRATE",
	OutTemp       => PPCS0PLBREARBITRATE_OUT,
	Paths         => (0 => (CPMPPCS0PLBCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS0PLBSSIZE(0),
	GlitchData    => PPCS0PLBSSIZE0_GlitchData,
	OutSignalName => "PPCS0PLBSSIZE(0)",
	OutTemp       => PPCS0PLBSSIZE_OUT(0),
	Paths         => (0 => (CPMPPCS0PLBCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS0PLBSSIZE(1),
	GlitchData    => PPCS0PLBSSIZE1_GlitchData,
	OutSignalName => "PPCS0PLBSSIZE(1)",
	OutTemp       => PPCS0PLBSSIZE_OUT(1),
	Paths         => (0 => (CPMPPCS0PLBCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS0PLBWAIT,
	GlitchData    => PPCS0PLBWAIT_GlitchData,
	OutSignalName => "PPCS0PLBWAIT",
	OutTemp       => PPCS0PLBWAIT_OUT,
	Paths         => (0 => (CPMPPCS0PLBCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS0PLBWRBTERM,
	GlitchData    => PPCS0PLBWRBTERM_GlitchData,
	OutSignalName => "PPCS0PLBWRBTERM",
	OutTemp       => PPCS0PLBWRBTERM_OUT,
	Paths         => (0 => (CPMPPCS0PLBCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS0PLBWRCOMP,
	GlitchData    => PPCS0PLBWRCOMP_GlitchData,
	OutSignalName => "PPCS0PLBWRCOMP",
	OutTemp       => PPCS0PLBWRCOMP_OUT,
	Paths         => (0 => (CPMPPCS0PLBCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS0PLBWRDACK,
	GlitchData    => PPCS0PLBWRDACK_GlitchData,
	OutSignalName => "PPCS0PLBWRDACK",
	OutTemp       => PPCS0PLBWRDACK_OUT,
	Paths         => (0 => (CPMPPCS0PLBCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS1PLBADDRACK,
	GlitchData    => PPCS1PLBADDRACK_GlitchData,
	OutSignalName => "PPCS1PLBADDRACK",
	OutTemp       => PPCS1PLBADDRACK_OUT,
	Paths         => (0 => (CPMPPCS1PLBCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS1PLBMBUSY(0),
	GlitchData    => PPCS1PLBMBUSY0_GlitchData,
	OutSignalName => "PPCS1PLBMBUSY(0)",
	OutTemp       => PPCS1PLBMBUSY_OUT(0),
	Paths         => (0 => (CPMPPCS1PLBCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS1PLBMBUSY(1),
	GlitchData    => PPCS1PLBMBUSY1_GlitchData,
	OutSignalName => "PPCS1PLBMBUSY(1)",
	OutTemp       => PPCS1PLBMBUSY_OUT(1),
	Paths         => (0 => (CPMPPCS1PLBCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS1PLBMBUSY(2),
	GlitchData    => PPCS1PLBMBUSY2_GlitchData,
	OutSignalName => "PPCS1PLBMBUSY(2)",
	OutTemp       => PPCS1PLBMBUSY_OUT(2),
	Paths         => (0 => (CPMPPCS1PLBCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS1PLBMBUSY(3),
	GlitchData    => PPCS1PLBMBUSY3_GlitchData,
	OutSignalName => "PPCS1PLBMBUSY(3)",
	OutTemp       => PPCS1PLBMBUSY_OUT(3),
	Paths         => (0 => (CPMPPCS1PLBCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS1PLBMIRQ(0),
	GlitchData    => PPCS1PLBMIRQ0_GlitchData,
	OutSignalName => "PPCS1PLBMIRQ(0)",
	OutTemp       => PPCS1PLBMIRQ_OUT(0),
	Paths         => (0 => (CPMPPCS1PLBCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS1PLBMIRQ(1),
	GlitchData    => PPCS1PLBMIRQ1_GlitchData,
	OutSignalName => "PPCS1PLBMIRQ(1)",
	OutTemp       => PPCS1PLBMIRQ_OUT(1),
	Paths         => (0 => (CPMPPCS1PLBCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS1PLBMIRQ(2),
	GlitchData    => PPCS1PLBMIRQ2_GlitchData,
	OutSignalName => "PPCS1PLBMIRQ(2)",
	OutTemp       => PPCS1PLBMIRQ_OUT(2),
	Paths         => (0 => (CPMPPCS1PLBCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS1PLBMIRQ(3),
	GlitchData    => PPCS1PLBMIRQ3_GlitchData,
	OutSignalName => "PPCS1PLBMIRQ(3)",
	OutTemp       => PPCS1PLBMIRQ_OUT(3),
	Paths         => (0 => (CPMPPCS1PLBCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS1PLBMRDERR(0),
	GlitchData    => PPCS1PLBMRDERR0_GlitchData,
	OutSignalName => "PPCS1PLBMRDERR(0)",
	OutTemp       => PPCS1PLBMRDERR_OUT(0),
	Paths         => (0 => (CPMPPCS1PLBCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS1PLBMRDERR(1),
	GlitchData    => PPCS1PLBMRDERR1_GlitchData,
	OutSignalName => "PPCS1PLBMRDERR(1)",
	OutTemp       => PPCS1PLBMRDERR_OUT(1),
	Paths         => (0 => (CPMPPCS1PLBCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS1PLBMRDERR(2),
	GlitchData    => PPCS1PLBMRDERR2_GlitchData,
	OutSignalName => "PPCS1PLBMRDERR(2)",
	OutTemp       => PPCS1PLBMRDERR_OUT(2),
	Paths         => (0 => (CPMPPCS1PLBCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS1PLBMRDERR(3),
	GlitchData    => PPCS1PLBMRDERR3_GlitchData,
	OutSignalName => "PPCS1PLBMRDERR(3)",
	OutTemp       => PPCS1PLBMRDERR_OUT(3),
	Paths         => (0 => (CPMPPCS1PLBCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS1PLBMWRERR(0),
	GlitchData    => PPCS1PLBMWRERR0_GlitchData,
	OutSignalName => "PPCS1PLBMWRERR(0)",
	OutTemp       => PPCS1PLBMWRERR_OUT(0),
	Paths         => (0 => (CPMPPCS1PLBCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS1PLBMWRERR(1),
	GlitchData    => PPCS1PLBMWRERR1_GlitchData,
	OutSignalName => "PPCS1PLBMWRERR(1)",
	OutTemp       => PPCS1PLBMWRERR_OUT(1),
	Paths         => (0 => (CPMPPCS1PLBCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS1PLBMWRERR(2),
	GlitchData    => PPCS1PLBMWRERR2_GlitchData,
	OutSignalName => "PPCS1PLBMWRERR(2)",
	OutTemp       => PPCS1PLBMWRERR_OUT(2),
	Paths         => (0 => (CPMPPCS1PLBCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS1PLBMWRERR(3),
	GlitchData    => PPCS1PLBMWRERR3_GlitchData,
	OutSignalName => "PPCS1PLBMWRERR(3)",
	OutTemp       => PPCS1PLBMWRERR_OUT(3),
	Paths         => (0 => (CPMPPCS1PLBCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS1PLBRDBTERM,
	GlitchData    => PPCS1PLBRDBTERM_GlitchData,
	OutSignalName => "PPCS1PLBRDBTERM",
	OutTemp       => PPCS1PLBRDBTERM_OUT,
	Paths         => (0 => (CPMPPCS1PLBCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS1PLBRDCOMP,
	GlitchData    => PPCS1PLBRDCOMP_GlitchData,
	OutSignalName => "PPCS1PLBRDCOMP",
	OutTemp       => PPCS1PLBRDCOMP_OUT,
	Paths         => (0 => (CPMPPCS1PLBCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS1PLBRDDACK,
	GlitchData    => PPCS1PLBRDDACK_GlitchData,
	OutSignalName => "PPCS1PLBRDDACK",
	OutTemp       => PPCS1PLBRDDACK_OUT,
	Paths         => (0 => (CPMPPCS1PLBCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS1PLBRDDBUS(0),
	GlitchData    => PPCS1PLBRDDBUS0_GlitchData,
	OutSignalName => "PPCS1PLBRDDBUS(0)",
	OutTemp       => PPCS1PLBRDDBUS_OUT(0),
	Paths         => (0 => (CPMPPCS1PLBCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS1PLBRDDBUS(1),
	GlitchData    => PPCS1PLBRDDBUS1_GlitchData,
	OutSignalName => "PPCS1PLBRDDBUS(1)",
	OutTemp       => PPCS1PLBRDDBUS_OUT(1),
	Paths         => (0 => (CPMPPCS1PLBCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS1PLBRDDBUS(2),
	GlitchData    => PPCS1PLBRDDBUS2_GlitchData,
	OutSignalName => "PPCS1PLBRDDBUS(2)",
	OutTemp       => PPCS1PLBRDDBUS_OUT(2),
	Paths         => (0 => (CPMPPCS1PLBCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS1PLBRDDBUS(3),
	GlitchData    => PPCS1PLBRDDBUS3_GlitchData,
	OutSignalName => "PPCS1PLBRDDBUS(3)",
	OutTemp       => PPCS1PLBRDDBUS_OUT(3),
	Paths         => (0 => (CPMPPCS1PLBCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS1PLBRDDBUS(4),
	GlitchData    => PPCS1PLBRDDBUS4_GlitchData,
	OutSignalName => "PPCS1PLBRDDBUS(4)",
	OutTemp       => PPCS1PLBRDDBUS_OUT(4),
	Paths         => (0 => (CPMPPCS1PLBCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS1PLBRDDBUS(5),
	GlitchData    => PPCS1PLBRDDBUS5_GlitchData,
	OutSignalName => "PPCS1PLBRDDBUS(5)",
	OutTemp       => PPCS1PLBRDDBUS_OUT(5),
	Paths         => (0 => (CPMPPCS1PLBCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS1PLBRDDBUS(6),
	GlitchData    => PPCS1PLBRDDBUS6_GlitchData,
	OutSignalName => "PPCS1PLBRDDBUS(6)",
	OutTemp       => PPCS1PLBRDDBUS_OUT(6),
	Paths         => (0 => (CPMPPCS1PLBCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS1PLBRDDBUS(7),
	GlitchData    => PPCS1PLBRDDBUS7_GlitchData,
	OutSignalName => "PPCS1PLBRDDBUS(7)",
	OutTemp       => PPCS1PLBRDDBUS_OUT(7),
	Paths         => (0 => (CPMPPCS1PLBCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS1PLBRDDBUS(8),
	GlitchData    => PPCS1PLBRDDBUS8_GlitchData,
	OutSignalName => "PPCS1PLBRDDBUS(8)",
	OutTemp       => PPCS1PLBRDDBUS_OUT(8),
	Paths         => (0 => (CPMPPCS1PLBCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS1PLBRDDBUS(9),
	GlitchData    => PPCS1PLBRDDBUS9_GlitchData,
	OutSignalName => "PPCS1PLBRDDBUS(9)",
	OutTemp       => PPCS1PLBRDDBUS_OUT(9),
	Paths         => (0 => (CPMPPCS1PLBCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS1PLBRDDBUS(10),
	GlitchData    => PPCS1PLBRDDBUS10_GlitchData,
	OutSignalName => "PPCS1PLBRDDBUS(10)",
	OutTemp       => PPCS1PLBRDDBUS_OUT(10),
	Paths         => (0 => (CPMPPCS1PLBCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS1PLBRDDBUS(11),
	GlitchData    => PPCS1PLBRDDBUS11_GlitchData,
	OutSignalName => "PPCS1PLBRDDBUS(11)",
	OutTemp       => PPCS1PLBRDDBUS_OUT(11),
	Paths         => (0 => (CPMPPCS1PLBCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS1PLBRDDBUS(12),
	GlitchData    => PPCS1PLBRDDBUS12_GlitchData,
	OutSignalName => "PPCS1PLBRDDBUS(12)",
	OutTemp       => PPCS1PLBRDDBUS_OUT(12),
	Paths         => (0 => (CPMPPCS1PLBCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS1PLBRDDBUS(13),
	GlitchData    => PPCS1PLBRDDBUS13_GlitchData,
	OutSignalName => "PPCS1PLBRDDBUS(13)",
	OutTemp       => PPCS1PLBRDDBUS_OUT(13),
	Paths         => (0 => (CPMPPCS1PLBCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS1PLBRDDBUS(14),
	GlitchData    => PPCS1PLBRDDBUS14_GlitchData,
	OutSignalName => "PPCS1PLBRDDBUS(14)",
	OutTemp       => PPCS1PLBRDDBUS_OUT(14),
	Paths         => (0 => (CPMPPCS1PLBCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS1PLBRDDBUS(15),
	GlitchData    => PPCS1PLBRDDBUS15_GlitchData,
	OutSignalName => "PPCS1PLBRDDBUS(15)",
	OutTemp       => PPCS1PLBRDDBUS_OUT(15),
	Paths         => (0 => (CPMPPCS1PLBCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS1PLBRDDBUS(16),
	GlitchData    => PPCS1PLBRDDBUS16_GlitchData,
	OutSignalName => "PPCS1PLBRDDBUS(16)",
	OutTemp       => PPCS1PLBRDDBUS_OUT(16),
	Paths         => (0 => (CPMPPCS1PLBCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS1PLBRDDBUS(17),
	GlitchData    => PPCS1PLBRDDBUS17_GlitchData,
	OutSignalName => "PPCS1PLBRDDBUS(17)",
	OutTemp       => PPCS1PLBRDDBUS_OUT(17),
	Paths         => (0 => (CPMPPCS1PLBCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS1PLBRDDBUS(18),
	GlitchData    => PPCS1PLBRDDBUS18_GlitchData,
	OutSignalName => "PPCS1PLBRDDBUS(18)",
	OutTemp       => PPCS1PLBRDDBUS_OUT(18),
	Paths         => (0 => (CPMPPCS1PLBCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS1PLBRDDBUS(19),
	GlitchData    => PPCS1PLBRDDBUS19_GlitchData,
	OutSignalName => "PPCS1PLBRDDBUS(19)",
	OutTemp       => PPCS1PLBRDDBUS_OUT(19),
	Paths         => (0 => (CPMPPCS1PLBCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS1PLBRDDBUS(20),
	GlitchData    => PPCS1PLBRDDBUS20_GlitchData,
	OutSignalName => "PPCS1PLBRDDBUS(20)",
	OutTemp       => PPCS1PLBRDDBUS_OUT(20),
	Paths         => (0 => (CPMPPCS1PLBCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS1PLBRDDBUS(21),
	GlitchData    => PPCS1PLBRDDBUS21_GlitchData,
	OutSignalName => "PPCS1PLBRDDBUS(21)",
	OutTemp       => PPCS1PLBRDDBUS_OUT(21),
	Paths         => (0 => (CPMPPCS1PLBCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS1PLBRDDBUS(22),
	GlitchData    => PPCS1PLBRDDBUS22_GlitchData,
	OutSignalName => "PPCS1PLBRDDBUS(22)",
	OutTemp       => PPCS1PLBRDDBUS_OUT(22),
	Paths         => (0 => (CPMPPCS1PLBCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS1PLBRDDBUS(23),
	GlitchData    => PPCS1PLBRDDBUS23_GlitchData,
	OutSignalName => "PPCS1PLBRDDBUS(23)",
	OutTemp       => PPCS1PLBRDDBUS_OUT(23),
	Paths         => (0 => (CPMPPCS1PLBCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS1PLBRDDBUS(24),
	GlitchData    => PPCS1PLBRDDBUS24_GlitchData,
	OutSignalName => "PPCS1PLBRDDBUS(24)",
	OutTemp       => PPCS1PLBRDDBUS_OUT(24),
	Paths         => (0 => (CPMPPCS1PLBCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS1PLBRDDBUS(25),
	GlitchData    => PPCS1PLBRDDBUS25_GlitchData,
	OutSignalName => "PPCS1PLBRDDBUS(25)",
	OutTemp       => PPCS1PLBRDDBUS_OUT(25),
	Paths         => (0 => (CPMPPCS1PLBCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS1PLBRDDBUS(26),
	GlitchData    => PPCS1PLBRDDBUS26_GlitchData,
	OutSignalName => "PPCS1PLBRDDBUS(26)",
	OutTemp       => PPCS1PLBRDDBUS_OUT(26),
	Paths         => (0 => (CPMPPCS1PLBCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS1PLBRDDBUS(27),
	GlitchData    => PPCS1PLBRDDBUS27_GlitchData,
	OutSignalName => "PPCS1PLBRDDBUS(27)",
	OutTemp       => PPCS1PLBRDDBUS_OUT(27),
	Paths         => (0 => (CPMPPCS1PLBCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS1PLBRDDBUS(28),
	GlitchData    => PPCS1PLBRDDBUS28_GlitchData,
	OutSignalName => "PPCS1PLBRDDBUS(28)",
	OutTemp       => PPCS1PLBRDDBUS_OUT(28),
	Paths         => (0 => (CPMPPCS1PLBCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS1PLBRDDBUS(29),
	GlitchData    => PPCS1PLBRDDBUS29_GlitchData,
	OutSignalName => "PPCS1PLBRDDBUS(29)",
	OutTemp       => PPCS1PLBRDDBUS_OUT(29),
	Paths         => (0 => (CPMPPCS1PLBCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS1PLBRDDBUS(30),
	GlitchData    => PPCS1PLBRDDBUS30_GlitchData,
	OutSignalName => "PPCS1PLBRDDBUS(30)",
	OutTemp       => PPCS1PLBRDDBUS_OUT(30),
	Paths         => (0 => (CPMPPCS1PLBCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS1PLBRDDBUS(31),
	GlitchData    => PPCS1PLBRDDBUS31_GlitchData,
	OutSignalName => "PPCS1PLBRDDBUS(31)",
	OutTemp       => PPCS1PLBRDDBUS_OUT(31),
	Paths         => (0 => (CPMPPCS1PLBCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS1PLBRDDBUS(32),
	GlitchData    => PPCS1PLBRDDBUS32_GlitchData,
	OutSignalName => "PPCS1PLBRDDBUS(32)",
	OutTemp       => PPCS1PLBRDDBUS_OUT(32),
	Paths         => (0 => (CPMPPCS1PLBCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS1PLBRDDBUS(33),
	GlitchData    => PPCS1PLBRDDBUS33_GlitchData,
	OutSignalName => "PPCS1PLBRDDBUS(33)",
	OutTemp       => PPCS1PLBRDDBUS_OUT(33),
	Paths         => (0 => (CPMPPCS1PLBCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS1PLBRDDBUS(34),
	GlitchData    => PPCS1PLBRDDBUS34_GlitchData,
	OutSignalName => "PPCS1PLBRDDBUS(34)",
	OutTemp       => PPCS1PLBRDDBUS_OUT(34),
	Paths         => (0 => (CPMPPCS1PLBCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS1PLBRDDBUS(35),
	GlitchData    => PPCS1PLBRDDBUS35_GlitchData,
	OutSignalName => "PPCS1PLBRDDBUS(35)",
	OutTemp       => PPCS1PLBRDDBUS_OUT(35),
	Paths         => (0 => (CPMPPCS1PLBCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS1PLBRDDBUS(36),
	GlitchData    => PPCS1PLBRDDBUS36_GlitchData,
	OutSignalName => "PPCS1PLBRDDBUS(36)",
	OutTemp       => PPCS1PLBRDDBUS_OUT(36),
	Paths         => (0 => (CPMPPCS1PLBCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS1PLBRDDBUS(37),
	GlitchData    => PPCS1PLBRDDBUS37_GlitchData,
	OutSignalName => "PPCS1PLBRDDBUS(37)",
	OutTemp       => PPCS1PLBRDDBUS_OUT(37),
	Paths         => (0 => (CPMPPCS1PLBCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS1PLBRDDBUS(38),
	GlitchData    => PPCS1PLBRDDBUS38_GlitchData,
	OutSignalName => "PPCS1PLBRDDBUS(38)",
	OutTemp       => PPCS1PLBRDDBUS_OUT(38),
	Paths         => (0 => (CPMPPCS1PLBCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS1PLBRDDBUS(39),
	GlitchData    => PPCS1PLBRDDBUS39_GlitchData,
	OutSignalName => "PPCS1PLBRDDBUS(39)",
	OutTemp       => PPCS1PLBRDDBUS_OUT(39),
	Paths         => (0 => (CPMPPCS1PLBCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS1PLBRDDBUS(40),
	GlitchData    => PPCS1PLBRDDBUS40_GlitchData,
	OutSignalName => "PPCS1PLBRDDBUS(40)",
	OutTemp       => PPCS1PLBRDDBUS_OUT(40),
	Paths         => (0 => (CPMPPCS1PLBCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS1PLBRDDBUS(41),
	GlitchData    => PPCS1PLBRDDBUS41_GlitchData,
	OutSignalName => "PPCS1PLBRDDBUS(41)",
	OutTemp       => PPCS1PLBRDDBUS_OUT(41),
	Paths         => (0 => (CPMPPCS1PLBCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS1PLBRDDBUS(42),
	GlitchData    => PPCS1PLBRDDBUS42_GlitchData,
	OutSignalName => "PPCS1PLBRDDBUS(42)",
	OutTemp       => PPCS1PLBRDDBUS_OUT(42),
	Paths         => (0 => (CPMPPCS1PLBCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS1PLBRDDBUS(43),
	GlitchData    => PPCS1PLBRDDBUS43_GlitchData,
	OutSignalName => "PPCS1PLBRDDBUS(43)",
	OutTemp       => PPCS1PLBRDDBUS_OUT(43),
	Paths         => (0 => (CPMPPCS1PLBCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS1PLBRDDBUS(44),
	GlitchData    => PPCS1PLBRDDBUS44_GlitchData,
	OutSignalName => "PPCS1PLBRDDBUS(44)",
	OutTemp       => PPCS1PLBRDDBUS_OUT(44),
	Paths         => (0 => (CPMPPCS1PLBCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS1PLBRDDBUS(45),
	GlitchData    => PPCS1PLBRDDBUS45_GlitchData,
	OutSignalName => "PPCS1PLBRDDBUS(45)",
	OutTemp       => PPCS1PLBRDDBUS_OUT(45),
	Paths         => (0 => (CPMPPCS1PLBCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS1PLBRDDBUS(46),
	GlitchData    => PPCS1PLBRDDBUS46_GlitchData,
	OutSignalName => "PPCS1PLBRDDBUS(46)",
	OutTemp       => PPCS1PLBRDDBUS_OUT(46),
	Paths         => (0 => (CPMPPCS1PLBCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS1PLBRDDBUS(47),
	GlitchData    => PPCS1PLBRDDBUS47_GlitchData,
	OutSignalName => "PPCS1PLBRDDBUS(47)",
	OutTemp       => PPCS1PLBRDDBUS_OUT(47),
	Paths         => (0 => (CPMPPCS1PLBCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS1PLBRDDBUS(48),
	GlitchData    => PPCS1PLBRDDBUS48_GlitchData,
	OutSignalName => "PPCS1PLBRDDBUS(48)",
	OutTemp       => PPCS1PLBRDDBUS_OUT(48),
	Paths         => (0 => (CPMPPCS1PLBCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS1PLBRDDBUS(49),
	GlitchData    => PPCS1PLBRDDBUS49_GlitchData,
	OutSignalName => "PPCS1PLBRDDBUS(49)",
	OutTemp       => PPCS1PLBRDDBUS_OUT(49),
	Paths         => (0 => (CPMPPCS1PLBCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS1PLBRDDBUS(50),
	GlitchData    => PPCS1PLBRDDBUS50_GlitchData,
	OutSignalName => "PPCS1PLBRDDBUS(50)",
	OutTemp       => PPCS1PLBRDDBUS_OUT(50),
	Paths         => (0 => (CPMPPCS1PLBCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS1PLBRDDBUS(51),
	GlitchData    => PPCS1PLBRDDBUS51_GlitchData,
	OutSignalName => "PPCS1PLBRDDBUS(51)",
	OutTemp       => PPCS1PLBRDDBUS_OUT(51),
	Paths         => (0 => (CPMPPCS1PLBCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS1PLBRDDBUS(52),
	GlitchData    => PPCS1PLBRDDBUS52_GlitchData,
	OutSignalName => "PPCS1PLBRDDBUS(52)",
	OutTemp       => PPCS1PLBRDDBUS_OUT(52),
	Paths         => (0 => (CPMPPCS1PLBCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS1PLBRDDBUS(53),
	GlitchData    => PPCS1PLBRDDBUS53_GlitchData,
	OutSignalName => "PPCS1PLBRDDBUS(53)",
	OutTemp       => PPCS1PLBRDDBUS_OUT(53),
	Paths         => (0 => (CPMPPCS1PLBCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS1PLBRDDBUS(54),
	GlitchData    => PPCS1PLBRDDBUS54_GlitchData,
	OutSignalName => "PPCS1PLBRDDBUS(54)",
	OutTemp       => PPCS1PLBRDDBUS_OUT(54),
	Paths         => (0 => (CPMPPCS1PLBCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS1PLBRDDBUS(55),
	GlitchData    => PPCS1PLBRDDBUS55_GlitchData,
	OutSignalName => "PPCS1PLBRDDBUS(55)",
	OutTemp       => PPCS1PLBRDDBUS_OUT(55),
	Paths         => (0 => (CPMPPCS1PLBCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS1PLBRDDBUS(56),
	GlitchData    => PPCS1PLBRDDBUS56_GlitchData,
	OutSignalName => "PPCS1PLBRDDBUS(56)",
	OutTemp       => PPCS1PLBRDDBUS_OUT(56),
	Paths         => (0 => (CPMPPCS1PLBCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS1PLBRDDBUS(57),
	GlitchData    => PPCS1PLBRDDBUS57_GlitchData,
	OutSignalName => "PPCS1PLBRDDBUS(57)",
	OutTemp       => PPCS1PLBRDDBUS_OUT(57),
	Paths         => (0 => (CPMPPCS1PLBCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS1PLBRDDBUS(58),
	GlitchData    => PPCS1PLBRDDBUS58_GlitchData,
	OutSignalName => "PPCS1PLBRDDBUS(58)",
	OutTemp       => PPCS1PLBRDDBUS_OUT(58),
	Paths         => (0 => (CPMPPCS1PLBCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS1PLBRDDBUS(59),
	GlitchData    => PPCS1PLBRDDBUS59_GlitchData,
	OutSignalName => "PPCS1PLBRDDBUS(59)",
	OutTemp       => PPCS1PLBRDDBUS_OUT(59),
	Paths         => (0 => (CPMPPCS1PLBCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS1PLBRDDBUS(60),
	GlitchData    => PPCS1PLBRDDBUS60_GlitchData,
	OutSignalName => "PPCS1PLBRDDBUS(60)",
	OutTemp       => PPCS1PLBRDDBUS_OUT(60),
	Paths         => (0 => (CPMPPCS1PLBCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS1PLBRDDBUS(61),
	GlitchData    => PPCS1PLBRDDBUS61_GlitchData,
	OutSignalName => "PPCS1PLBRDDBUS(61)",
	OutTemp       => PPCS1PLBRDDBUS_OUT(61),
	Paths         => (0 => (CPMPPCS1PLBCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS1PLBRDDBUS(62),
	GlitchData    => PPCS1PLBRDDBUS62_GlitchData,
	OutSignalName => "PPCS1PLBRDDBUS(62)",
	OutTemp       => PPCS1PLBRDDBUS_OUT(62),
	Paths         => (0 => (CPMPPCS1PLBCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS1PLBRDDBUS(63),
	GlitchData    => PPCS1PLBRDDBUS63_GlitchData,
	OutSignalName => "PPCS1PLBRDDBUS(63)",
	OutTemp       => PPCS1PLBRDDBUS_OUT(63),
	Paths         => (0 => (CPMPPCS1PLBCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS1PLBRDDBUS(64),
	GlitchData    => PPCS1PLBRDDBUS64_GlitchData,
	OutSignalName => "PPCS1PLBRDDBUS(64)",
	OutTemp       => PPCS1PLBRDDBUS_OUT(64),
	Paths         => (0 => (CPMPPCS1PLBCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS1PLBRDDBUS(65),
	GlitchData    => PPCS1PLBRDDBUS65_GlitchData,
	OutSignalName => "PPCS1PLBRDDBUS(65)",
	OutTemp       => PPCS1PLBRDDBUS_OUT(65),
	Paths         => (0 => (CPMPPCS1PLBCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS1PLBRDDBUS(66),
	GlitchData    => PPCS1PLBRDDBUS66_GlitchData,
	OutSignalName => "PPCS1PLBRDDBUS(66)",
	OutTemp       => PPCS1PLBRDDBUS_OUT(66),
	Paths         => (0 => (CPMPPCS1PLBCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS1PLBRDDBUS(67),
	GlitchData    => PPCS1PLBRDDBUS67_GlitchData,
	OutSignalName => "PPCS1PLBRDDBUS(67)",
	OutTemp       => PPCS1PLBRDDBUS_OUT(67),
	Paths         => (0 => (CPMPPCS1PLBCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS1PLBRDDBUS(68),
	GlitchData    => PPCS1PLBRDDBUS68_GlitchData,
	OutSignalName => "PPCS1PLBRDDBUS(68)",
	OutTemp       => PPCS1PLBRDDBUS_OUT(68),
	Paths         => (0 => (CPMPPCS1PLBCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS1PLBRDDBUS(69),
	GlitchData    => PPCS1PLBRDDBUS69_GlitchData,
	OutSignalName => "PPCS1PLBRDDBUS(69)",
	OutTemp       => PPCS1PLBRDDBUS_OUT(69),
	Paths         => (0 => (CPMPPCS1PLBCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS1PLBRDDBUS(70),
	GlitchData    => PPCS1PLBRDDBUS70_GlitchData,
	OutSignalName => "PPCS1PLBRDDBUS(70)",
	OutTemp       => PPCS1PLBRDDBUS_OUT(70),
	Paths         => (0 => (CPMPPCS1PLBCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS1PLBRDDBUS(71),
	GlitchData    => PPCS1PLBRDDBUS71_GlitchData,
	OutSignalName => "PPCS1PLBRDDBUS(71)",
	OutTemp       => PPCS1PLBRDDBUS_OUT(71),
	Paths         => (0 => (CPMPPCS1PLBCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS1PLBRDDBUS(72),
	GlitchData    => PPCS1PLBRDDBUS72_GlitchData,
	OutSignalName => "PPCS1PLBRDDBUS(72)",
	OutTemp       => PPCS1PLBRDDBUS_OUT(72),
	Paths         => (0 => (CPMPPCS1PLBCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS1PLBRDDBUS(73),
	GlitchData    => PPCS1PLBRDDBUS73_GlitchData,
	OutSignalName => "PPCS1PLBRDDBUS(73)",
	OutTemp       => PPCS1PLBRDDBUS_OUT(73),
	Paths         => (0 => (CPMPPCS1PLBCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS1PLBRDDBUS(74),
	GlitchData    => PPCS1PLBRDDBUS74_GlitchData,
	OutSignalName => "PPCS1PLBRDDBUS(74)",
	OutTemp       => PPCS1PLBRDDBUS_OUT(74),
	Paths         => (0 => (CPMPPCS1PLBCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS1PLBRDDBUS(75),
	GlitchData    => PPCS1PLBRDDBUS75_GlitchData,
	OutSignalName => "PPCS1PLBRDDBUS(75)",
	OutTemp       => PPCS1PLBRDDBUS_OUT(75),
	Paths         => (0 => (CPMPPCS1PLBCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS1PLBRDDBUS(76),
	GlitchData    => PPCS1PLBRDDBUS76_GlitchData,
	OutSignalName => "PPCS1PLBRDDBUS(76)",
	OutTemp       => PPCS1PLBRDDBUS_OUT(76),
	Paths         => (0 => (CPMPPCS1PLBCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS1PLBRDDBUS(77),
	GlitchData    => PPCS1PLBRDDBUS77_GlitchData,
	OutSignalName => "PPCS1PLBRDDBUS(77)",
	OutTemp       => PPCS1PLBRDDBUS_OUT(77),
	Paths         => (0 => (CPMPPCS1PLBCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS1PLBRDDBUS(78),
	GlitchData    => PPCS1PLBRDDBUS78_GlitchData,
	OutSignalName => "PPCS1PLBRDDBUS(78)",
	OutTemp       => PPCS1PLBRDDBUS_OUT(78),
	Paths         => (0 => (CPMPPCS1PLBCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS1PLBRDDBUS(79),
	GlitchData    => PPCS1PLBRDDBUS79_GlitchData,
	OutSignalName => "PPCS1PLBRDDBUS(79)",
	OutTemp       => PPCS1PLBRDDBUS_OUT(79),
	Paths         => (0 => (CPMPPCS1PLBCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS1PLBRDDBUS(80),
	GlitchData    => PPCS1PLBRDDBUS80_GlitchData,
	OutSignalName => "PPCS1PLBRDDBUS(80)",
	OutTemp       => PPCS1PLBRDDBUS_OUT(80),
	Paths         => (0 => (CPMPPCS1PLBCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS1PLBRDDBUS(81),
	GlitchData    => PPCS1PLBRDDBUS81_GlitchData,
	OutSignalName => "PPCS1PLBRDDBUS(81)",
	OutTemp       => PPCS1PLBRDDBUS_OUT(81),
	Paths         => (0 => (CPMPPCS1PLBCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS1PLBRDDBUS(82),
	GlitchData    => PPCS1PLBRDDBUS82_GlitchData,
	OutSignalName => "PPCS1PLBRDDBUS(82)",
	OutTemp       => PPCS1PLBRDDBUS_OUT(82),
	Paths         => (0 => (CPMPPCS1PLBCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS1PLBRDDBUS(83),
	GlitchData    => PPCS1PLBRDDBUS83_GlitchData,
	OutSignalName => "PPCS1PLBRDDBUS(83)",
	OutTemp       => PPCS1PLBRDDBUS_OUT(83),
	Paths         => (0 => (CPMPPCS1PLBCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS1PLBRDDBUS(84),
	GlitchData    => PPCS1PLBRDDBUS84_GlitchData,
	OutSignalName => "PPCS1PLBRDDBUS(84)",
	OutTemp       => PPCS1PLBRDDBUS_OUT(84),
	Paths         => (0 => (CPMPPCS1PLBCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS1PLBRDDBUS(85),
	GlitchData    => PPCS1PLBRDDBUS85_GlitchData,
	OutSignalName => "PPCS1PLBRDDBUS(85)",
	OutTemp       => PPCS1PLBRDDBUS_OUT(85),
	Paths         => (0 => (CPMPPCS1PLBCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS1PLBRDDBUS(86),
	GlitchData    => PPCS1PLBRDDBUS86_GlitchData,
	OutSignalName => "PPCS1PLBRDDBUS(86)",
	OutTemp       => PPCS1PLBRDDBUS_OUT(86),
	Paths         => (0 => (CPMPPCS1PLBCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS1PLBRDDBUS(87),
	GlitchData    => PPCS1PLBRDDBUS87_GlitchData,
	OutSignalName => "PPCS1PLBRDDBUS(87)",
	OutTemp       => PPCS1PLBRDDBUS_OUT(87),
	Paths         => (0 => (CPMPPCS1PLBCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS1PLBRDDBUS(88),
	GlitchData    => PPCS1PLBRDDBUS88_GlitchData,
	OutSignalName => "PPCS1PLBRDDBUS(88)",
	OutTemp       => PPCS1PLBRDDBUS_OUT(88),
	Paths         => (0 => (CPMPPCS1PLBCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS1PLBRDDBUS(89),
	GlitchData    => PPCS1PLBRDDBUS89_GlitchData,
	OutSignalName => "PPCS1PLBRDDBUS(89)",
	OutTemp       => PPCS1PLBRDDBUS_OUT(89),
	Paths         => (0 => (CPMPPCS1PLBCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS1PLBRDDBUS(90),
	GlitchData    => PPCS1PLBRDDBUS90_GlitchData,
	OutSignalName => "PPCS1PLBRDDBUS(90)",
	OutTemp       => PPCS1PLBRDDBUS_OUT(90),
	Paths         => (0 => (CPMPPCS1PLBCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS1PLBRDDBUS(91),
	GlitchData    => PPCS1PLBRDDBUS91_GlitchData,
	OutSignalName => "PPCS1PLBRDDBUS(91)",
	OutTemp       => PPCS1PLBRDDBUS_OUT(91),
	Paths         => (0 => (CPMPPCS1PLBCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS1PLBRDDBUS(92),
	GlitchData    => PPCS1PLBRDDBUS92_GlitchData,
	OutSignalName => "PPCS1PLBRDDBUS(92)",
	OutTemp       => PPCS1PLBRDDBUS_OUT(92),
	Paths         => (0 => (CPMPPCS1PLBCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS1PLBRDDBUS(93),
	GlitchData    => PPCS1PLBRDDBUS93_GlitchData,
	OutSignalName => "PPCS1PLBRDDBUS(93)",
	OutTemp       => PPCS1PLBRDDBUS_OUT(93),
	Paths         => (0 => (CPMPPCS1PLBCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS1PLBRDDBUS(94),
	GlitchData    => PPCS1PLBRDDBUS94_GlitchData,
	OutSignalName => "PPCS1PLBRDDBUS(94)",
	OutTemp       => PPCS1PLBRDDBUS_OUT(94),
	Paths         => (0 => (CPMPPCS1PLBCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS1PLBRDDBUS(95),
	GlitchData    => PPCS1PLBRDDBUS95_GlitchData,
	OutSignalName => "PPCS1PLBRDDBUS(95)",
	OutTemp       => PPCS1PLBRDDBUS_OUT(95),
	Paths         => (0 => (CPMPPCS1PLBCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS1PLBRDDBUS(96),
	GlitchData    => PPCS1PLBRDDBUS96_GlitchData,
	OutSignalName => "PPCS1PLBRDDBUS(96)",
	OutTemp       => PPCS1PLBRDDBUS_OUT(96),
	Paths         => (0 => (CPMPPCS1PLBCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS1PLBRDDBUS(97),
	GlitchData    => PPCS1PLBRDDBUS97_GlitchData,
	OutSignalName => "PPCS1PLBRDDBUS(97)",
	OutTemp       => PPCS1PLBRDDBUS_OUT(97),
	Paths         => (0 => (CPMPPCS1PLBCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS1PLBRDDBUS(98),
	GlitchData    => PPCS1PLBRDDBUS98_GlitchData,
	OutSignalName => "PPCS1PLBRDDBUS(98)",
	OutTemp       => PPCS1PLBRDDBUS_OUT(98),
	Paths         => (0 => (CPMPPCS1PLBCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS1PLBRDDBUS(99),
	GlitchData    => PPCS1PLBRDDBUS99_GlitchData,
	OutSignalName => "PPCS1PLBRDDBUS(99)",
	OutTemp       => PPCS1PLBRDDBUS_OUT(99),
	Paths         => (0 => (CPMPPCS1PLBCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS1PLBRDDBUS(100),
	GlitchData    => PPCS1PLBRDDBUS100_GlitchData,
	OutSignalName => "PPCS1PLBRDDBUS(100)",
	OutTemp       => PPCS1PLBRDDBUS_OUT(100),
	Paths         => (0 => (CPMPPCS1PLBCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS1PLBRDDBUS(101),
	GlitchData    => PPCS1PLBRDDBUS101_GlitchData,
	OutSignalName => "PPCS1PLBRDDBUS(101)",
	OutTemp       => PPCS1PLBRDDBUS_OUT(101),
	Paths         => (0 => (CPMPPCS1PLBCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS1PLBRDDBUS(102),
	GlitchData    => PPCS1PLBRDDBUS102_GlitchData,
	OutSignalName => "PPCS1PLBRDDBUS(102)",
	OutTemp       => PPCS1PLBRDDBUS_OUT(102),
	Paths         => (0 => (CPMPPCS1PLBCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS1PLBRDDBUS(103),
	GlitchData    => PPCS1PLBRDDBUS103_GlitchData,
	OutSignalName => "PPCS1PLBRDDBUS(103)",
	OutTemp       => PPCS1PLBRDDBUS_OUT(103),
	Paths         => (0 => (CPMPPCS1PLBCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS1PLBRDDBUS(104),
	GlitchData    => PPCS1PLBRDDBUS104_GlitchData,
	OutSignalName => "PPCS1PLBRDDBUS(104)",
	OutTemp       => PPCS1PLBRDDBUS_OUT(104),
	Paths         => (0 => (CPMPPCS1PLBCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS1PLBRDDBUS(105),
	GlitchData    => PPCS1PLBRDDBUS105_GlitchData,
	OutSignalName => "PPCS1PLBRDDBUS(105)",
	OutTemp       => PPCS1PLBRDDBUS_OUT(105),
	Paths         => (0 => (CPMPPCS1PLBCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS1PLBRDDBUS(106),
	GlitchData    => PPCS1PLBRDDBUS106_GlitchData,
	OutSignalName => "PPCS1PLBRDDBUS(106)",
	OutTemp       => PPCS1PLBRDDBUS_OUT(106),
	Paths         => (0 => (CPMPPCS1PLBCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS1PLBRDDBUS(107),
	GlitchData    => PPCS1PLBRDDBUS107_GlitchData,
	OutSignalName => "PPCS1PLBRDDBUS(107)",
	OutTemp       => PPCS1PLBRDDBUS_OUT(107),
	Paths         => (0 => (CPMPPCS1PLBCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS1PLBRDDBUS(108),
	GlitchData    => PPCS1PLBRDDBUS108_GlitchData,
	OutSignalName => "PPCS1PLBRDDBUS(108)",
	OutTemp       => PPCS1PLBRDDBUS_OUT(108),
	Paths         => (0 => (CPMPPCS1PLBCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS1PLBRDDBUS(109),
	GlitchData    => PPCS1PLBRDDBUS109_GlitchData,
	OutSignalName => "PPCS1PLBRDDBUS(109)",
	OutTemp       => PPCS1PLBRDDBUS_OUT(109),
	Paths         => (0 => (CPMPPCS1PLBCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS1PLBRDDBUS(110),
	GlitchData    => PPCS1PLBRDDBUS110_GlitchData,
	OutSignalName => "PPCS1PLBRDDBUS(110)",
	OutTemp       => PPCS1PLBRDDBUS_OUT(110),
	Paths         => (0 => (CPMPPCS1PLBCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS1PLBRDDBUS(111),
	GlitchData    => PPCS1PLBRDDBUS111_GlitchData,
	OutSignalName => "PPCS1PLBRDDBUS(111)",
	OutTemp       => PPCS1PLBRDDBUS_OUT(111),
	Paths         => (0 => (CPMPPCS1PLBCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS1PLBRDDBUS(112),
	GlitchData    => PPCS1PLBRDDBUS112_GlitchData,
	OutSignalName => "PPCS1PLBRDDBUS(112)",
	OutTemp       => PPCS1PLBRDDBUS_OUT(112),
	Paths         => (0 => (CPMPPCS1PLBCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS1PLBRDDBUS(113),
	GlitchData    => PPCS1PLBRDDBUS113_GlitchData,
	OutSignalName => "PPCS1PLBRDDBUS(113)",
	OutTemp       => PPCS1PLBRDDBUS_OUT(113),
	Paths         => (0 => (CPMPPCS1PLBCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS1PLBRDDBUS(114),
	GlitchData    => PPCS1PLBRDDBUS114_GlitchData,
	OutSignalName => "PPCS1PLBRDDBUS(114)",
	OutTemp       => PPCS1PLBRDDBUS_OUT(114),
	Paths         => (0 => (CPMPPCS1PLBCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS1PLBRDDBUS(115),
	GlitchData    => PPCS1PLBRDDBUS115_GlitchData,
	OutSignalName => "PPCS1PLBRDDBUS(115)",
	OutTemp       => PPCS1PLBRDDBUS_OUT(115),
	Paths         => (0 => (CPMPPCS1PLBCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS1PLBRDDBUS(116),
	GlitchData    => PPCS1PLBRDDBUS116_GlitchData,
	OutSignalName => "PPCS1PLBRDDBUS(116)",
	OutTemp       => PPCS1PLBRDDBUS_OUT(116),
	Paths         => (0 => (CPMPPCS1PLBCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS1PLBRDDBUS(117),
	GlitchData    => PPCS1PLBRDDBUS117_GlitchData,
	OutSignalName => "PPCS1PLBRDDBUS(117)",
	OutTemp       => PPCS1PLBRDDBUS_OUT(117),
	Paths         => (0 => (CPMPPCS1PLBCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS1PLBRDDBUS(118),
	GlitchData    => PPCS1PLBRDDBUS118_GlitchData,
	OutSignalName => "PPCS1PLBRDDBUS(118)",
	OutTemp       => PPCS1PLBRDDBUS_OUT(118),
	Paths         => (0 => (CPMPPCS1PLBCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS1PLBRDDBUS(119),
	GlitchData    => PPCS1PLBRDDBUS119_GlitchData,
	OutSignalName => "PPCS1PLBRDDBUS(119)",
	OutTemp       => PPCS1PLBRDDBUS_OUT(119),
	Paths         => (0 => (CPMPPCS1PLBCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS1PLBRDDBUS(120),
	GlitchData    => PPCS1PLBRDDBUS120_GlitchData,
	OutSignalName => "PPCS1PLBRDDBUS(120)",
	OutTemp       => PPCS1PLBRDDBUS_OUT(120),
	Paths         => (0 => (CPMPPCS1PLBCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS1PLBRDDBUS(121),
	GlitchData    => PPCS1PLBRDDBUS121_GlitchData,
	OutSignalName => "PPCS1PLBRDDBUS(121)",
	OutTemp       => PPCS1PLBRDDBUS_OUT(121),
	Paths         => (0 => (CPMPPCS1PLBCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS1PLBRDDBUS(122),
	GlitchData    => PPCS1PLBRDDBUS122_GlitchData,
	OutSignalName => "PPCS1PLBRDDBUS(122)",
	OutTemp       => PPCS1PLBRDDBUS_OUT(122),
	Paths         => (0 => (CPMPPCS1PLBCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS1PLBRDDBUS(123),
	GlitchData    => PPCS1PLBRDDBUS123_GlitchData,
	OutSignalName => "PPCS1PLBRDDBUS(123)",
	OutTemp       => PPCS1PLBRDDBUS_OUT(123),
	Paths         => (0 => (CPMPPCS1PLBCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS1PLBRDDBUS(124),
	GlitchData    => PPCS1PLBRDDBUS124_GlitchData,
	OutSignalName => "PPCS1PLBRDDBUS(124)",
	OutTemp       => PPCS1PLBRDDBUS_OUT(124),
	Paths         => (0 => (CPMPPCS1PLBCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS1PLBRDDBUS(125),
	GlitchData    => PPCS1PLBRDDBUS125_GlitchData,
	OutSignalName => "PPCS1PLBRDDBUS(125)",
	OutTemp       => PPCS1PLBRDDBUS_OUT(125),
	Paths         => (0 => (CPMPPCS1PLBCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS1PLBRDDBUS(126),
	GlitchData    => PPCS1PLBRDDBUS126_GlitchData,
	OutSignalName => "PPCS1PLBRDDBUS(126)",
	OutTemp       => PPCS1PLBRDDBUS_OUT(126),
	Paths         => (0 => (CPMPPCS1PLBCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS1PLBRDDBUS(127),
	GlitchData    => PPCS1PLBRDDBUS127_GlitchData,
	OutSignalName => "PPCS1PLBRDDBUS(127)",
	OutTemp       => PPCS1PLBRDDBUS_OUT(127),
	Paths         => (0 => (CPMPPCS1PLBCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS1PLBRDWDADDR(0),
	GlitchData    => PPCS1PLBRDWDADDR0_GlitchData,
	OutSignalName => "PPCS1PLBRDWDADDR(0)",
	OutTemp       => PPCS1PLBRDWDADDR_OUT(0),
	Paths         => (0 => (CPMPPCS1PLBCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS1PLBRDWDADDR(1),
	GlitchData    => PPCS1PLBRDWDADDR1_GlitchData,
	OutSignalName => "PPCS1PLBRDWDADDR(1)",
	OutTemp       => PPCS1PLBRDWDADDR_OUT(1),
	Paths         => (0 => (CPMPPCS1PLBCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS1PLBRDWDADDR(2),
	GlitchData    => PPCS1PLBRDWDADDR2_GlitchData,
	OutSignalName => "PPCS1PLBRDWDADDR(2)",
	OutTemp       => PPCS1PLBRDWDADDR_OUT(2),
	Paths         => (0 => (CPMPPCS1PLBCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS1PLBRDWDADDR(3),
	GlitchData    => PPCS1PLBRDWDADDR3_GlitchData,
	OutSignalName => "PPCS1PLBRDWDADDR(3)",
	OutTemp       => PPCS1PLBRDWDADDR_OUT(3),
	Paths         => (0 => (CPMPPCS1PLBCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS1PLBREARBITRATE,
	GlitchData    => PPCS1PLBREARBITRATE_GlitchData,
	OutSignalName => "PPCS1PLBREARBITRATE",
	OutTemp       => PPCS1PLBREARBITRATE_OUT,
	Paths         => (0 => (CPMPPCS1PLBCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS1PLBSSIZE(0),
	GlitchData    => PPCS1PLBSSIZE0_GlitchData,
	OutSignalName => "PPCS1PLBSSIZE(0)",
	OutTemp       => PPCS1PLBSSIZE_OUT(0),
	Paths         => (0 => (CPMPPCS1PLBCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS1PLBSSIZE(1),
	GlitchData    => PPCS1PLBSSIZE1_GlitchData,
	OutSignalName => "PPCS1PLBSSIZE(1)",
	OutTemp       => PPCS1PLBSSIZE_OUT(1),
	Paths         => (0 => (CPMPPCS1PLBCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS1PLBWAIT,
	GlitchData    => PPCS1PLBWAIT_GlitchData,
	OutSignalName => "PPCS1PLBWAIT",
	OutTemp       => PPCS1PLBWAIT_OUT,
	Paths         => (0 => (CPMPPCS1PLBCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS1PLBWRBTERM,
	GlitchData    => PPCS1PLBWRBTERM_GlitchData,
	OutSignalName => "PPCS1PLBWRBTERM",
	OutTemp       => PPCS1PLBWRBTERM_OUT,
	Paths         => (0 => (CPMPPCS1PLBCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS1PLBWRCOMP,
	GlitchData    => PPCS1PLBWRCOMP_GlitchData,
	OutSignalName => "PPCS1PLBWRCOMP",
	OutTemp       => PPCS1PLBWRCOMP_OUT,
	Paths         => (0 => (CPMPPCS1PLBCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS1PLBWRDACK,
	GlitchData    => PPCS1PLBWRDACK_GlitchData,
	OutSignalName => "PPCS1PLBWRDACK",
	OutTemp       => PPCS1PLBWRDACK_OUT,
	Paths         => (0 => (CPMPPCS1PLBCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => APUFCMDECFPUOP,
	GlitchData    => APUFCMDECFPUOP_GlitchData,
	OutSignalName => "APUFCMDECFPUOP",
	OutTemp       => APUFCMDECFPUOP_OUT,
	Paths         => (0 => (CPMFCMCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => APUFCMDECLDSTXFERSIZE(0),
	GlitchData    => APUFCMDECLDSTXFERSIZE0_GlitchData,
	OutSignalName => "APUFCMDECLDSTXFERSIZE(0)",
	OutTemp       => APUFCMDECLDSTXFERSIZE_OUT(0),
	Paths         => (0 => (CPMFCMCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => APUFCMDECLDSTXFERSIZE(1),
	GlitchData    => APUFCMDECLDSTXFERSIZE1_GlitchData,
	OutSignalName => "APUFCMDECLDSTXFERSIZE(1)",
	OutTemp       => APUFCMDECLDSTXFERSIZE_OUT(1),
	Paths         => (0 => (CPMFCMCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => APUFCMDECLDSTXFERSIZE(2),
	GlitchData    => APUFCMDECLDSTXFERSIZE2_GlitchData,
	OutSignalName => "APUFCMDECLDSTXFERSIZE(2)",
	OutTemp       => APUFCMDECLDSTXFERSIZE_OUT(2),
	Paths         => (0 => (CPMFCMCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => APUFCMDECLOAD,
	GlitchData    => APUFCMDECLOAD_GlitchData,
	OutSignalName => "APUFCMDECLOAD",
	OutTemp       => APUFCMDECLOAD_OUT,
	Paths         => (0 => (CPMFCMCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => APUFCMDECNONAUTON,
	GlitchData    => APUFCMDECNONAUTON_GlitchData,
	OutSignalName => "APUFCMDECNONAUTON",
	OutTemp       => APUFCMDECNONAUTON_OUT,
	Paths         => (0 => (CPMFCMCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => APUFCMDECSTORE,
	GlitchData    => APUFCMDECSTORE_GlitchData,
	OutSignalName => "APUFCMDECSTORE",
	OutTemp       => APUFCMDECSTORE_OUT,
	Paths         => (0 => (CPMFCMCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => APUFCMDECUDI(0),
	GlitchData    => APUFCMDECUDI0_GlitchData,
	OutSignalName => "APUFCMDECUDI(0)",
	OutTemp       => APUFCMDECUDI_OUT(0),
	Paths         => (0 => (CPMFCMCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => APUFCMDECUDI(1),
	GlitchData    => APUFCMDECUDI1_GlitchData,
	OutSignalName => "APUFCMDECUDI(1)",
	OutTemp       => APUFCMDECUDI_OUT(1),
	Paths         => (0 => (CPMFCMCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => APUFCMDECUDI(2),
	GlitchData    => APUFCMDECUDI2_GlitchData,
	OutSignalName => "APUFCMDECUDI(2)",
	OutTemp       => APUFCMDECUDI_OUT(2),
	Paths         => (0 => (CPMFCMCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => APUFCMDECUDI(3),
	GlitchData    => APUFCMDECUDI3_GlitchData,
	OutSignalName => "APUFCMDECUDI(3)",
	OutTemp       => APUFCMDECUDI_OUT(3),
	Paths         => (0 => (CPMFCMCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => APUFCMDECUDIVALID,
	GlitchData    => APUFCMDECUDIVALID_GlitchData,
	OutSignalName => "APUFCMDECUDIVALID",
	OutTemp       => APUFCMDECUDIVALID_OUT,
	Paths         => (0 => (CPMFCMCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => APUFCMENDIAN,
	GlitchData    => APUFCMENDIAN_GlitchData,
	OutSignalName => "APUFCMENDIAN",
	OutTemp       => APUFCMENDIAN_OUT,
	Paths         => (0 => (CPMFCMCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => APUFCMFLUSH,
	GlitchData    => APUFCMFLUSH_GlitchData,
	OutSignalName => "APUFCMFLUSH",
	OutTemp       => APUFCMFLUSH_OUT,
	Paths         => (0 => (CPMFCMCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => APUFCMINSTRUCTION(0),
	GlitchData    => APUFCMINSTRUCTION0_GlitchData,
	OutSignalName => "APUFCMINSTRUCTION(0)",
	OutTemp       => APUFCMINSTRUCTION_OUT(0),
	Paths         => (0 => (CPMFCMCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => APUFCMINSTRUCTION(1),
	GlitchData    => APUFCMINSTRUCTION1_GlitchData,
	OutSignalName => "APUFCMINSTRUCTION(1)",
	OutTemp       => APUFCMINSTRUCTION_OUT(1),
	Paths         => (0 => (CPMFCMCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => APUFCMINSTRUCTION(2),
	GlitchData    => APUFCMINSTRUCTION2_GlitchData,
	OutSignalName => "APUFCMINSTRUCTION(2)",
	OutTemp       => APUFCMINSTRUCTION_OUT(2),
	Paths         => (0 => (CPMFCMCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => APUFCMINSTRUCTION(3),
	GlitchData    => APUFCMINSTRUCTION3_GlitchData,
	OutSignalName => "APUFCMINSTRUCTION(3)",
	OutTemp       => APUFCMINSTRUCTION_OUT(3),
	Paths         => (0 => (CPMFCMCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => APUFCMINSTRUCTION(4),
	GlitchData    => APUFCMINSTRUCTION4_GlitchData,
	OutSignalName => "APUFCMINSTRUCTION(4)",
	OutTemp       => APUFCMINSTRUCTION_OUT(4),
	Paths         => (0 => (CPMFCMCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => APUFCMINSTRUCTION(5),
	GlitchData    => APUFCMINSTRUCTION5_GlitchData,
	OutSignalName => "APUFCMINSTRUCTION(5)",
	OutTemp       => APUFCMINSTRUCTION_OUT(5),
	Paths         => (0 => (CPMFCMCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => APUFCMINSTRUCTION(6),
	GlitchData    => APUFCMINSTRUCTION6_GlitchData,
	OutSignalName => "APUFCMINSTRUCTION(6)",
	OutTemp       => APUFCMINSTRUCTION_OUT(6),
	Paths         => (0 => (CPMFCMCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => APUFCMINSTRUCTION(7),
	GlitchData    => APUFCMINSTRUCTION7_GlitchData,
	OutSignalName => "APUFCMINSTRUCTION(7)",
	OutTemp       => APUFCMINSTRUCTION_OUT(7),
	Paths         => (0 => (CPMFCMCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => APUFCMINSTRUCTION(8),
	GlitchData    => APUFCMINSTRUCTION8_GlitchData,
	OutSignalName => "APUFCMINSTRUCTION(8)",
	OutTemp       => APUFCMINSTRUCTION_OUT(8),
	Paths         => (0 => (CPMFCMCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => APUFCMINSTRUCTION(9),
	GlitchData    => APUFCMINSTRUCTION9_GlitchData,
	OutSignalName => "APUFCMINSTRUCTION(9)",
	OutTemp       => APUFCMINSTRUCTION_OUT(9),
	Paths         => (0 => (CPMFCMCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => APUFCMINSTRUCTION(10),
	GlitchData    => APUFCMINSTRUCTION10_GlitchData,
	OutSignalName => "APUFCMINSTRUCTION(10)",
	OutTemp       => APUFCMINSTRUCTION_OUT(10),
	Paths         => (0 => (CPMFCMCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => APUFCMINSTRUCTION(11),
	GlitchData    => APUFCMINSTRUCTION11_GlitchData,
	OutSignalName => "APUFCMINSTRUCTION(11)",
	OutTemp       => APUFCMINSTRUCTION_OUT(11),
	Paths         => (0 => (CPMFCMCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => APUFCMINSTRUCTION(12),
	GlitchData    => APUFCMINSTRUCTION12_GlitchData,
	OutSignalName => "APUFCMINSTRUCTION(12)",
	OutTemp       => APUFCMINSTRUCTION_OUT(12),
	Paths         => (0 => (CPMFCMCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => APUFCMINSTRUCTION(13),
	GlitchData    => APUFCMINSTRUCTION13_GlitchData,
	OutSignalName => "APUFCMINSTRUCTION(13)",
	OutTemp       => APUFCMINSTRUCTION_OUT(13),
	Paths         => (0 => (CPMFCMCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => APUFCMINSTRUCTION(14),
	GlitchData    => APUFCMINSTRUCTION14_GlitchData,
	OutSignalName => "APUFCMINSTRUCTION(14)",
	OutTemp       => APUFCMINSTRUCTION_OUT(14),
	Paths         => (0 => (CPMFCMCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => APUFCMINSTRUCTION(15),
	GlitchData    => APUFCMINSTRUCTION15_GlitchData,
	OutSignalName => "APUFCMINSTRUCTION(15)",
	OutTemp       => APUFCMINSTRUCTION_OUT(15),
	Paths         => (0 => (CPMFCMCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => APUFCMINSTRUCTION(16),
	GlitchData    => APUFCMINSTRUCTION16_GlitchData,
	OutSignalName => "APUFCMINSTRUCTION(16)",
	OutTemp       => APUFCMINSTRUCTION_OUT(16),
	Paths         => (0 => (CPMFCMCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => APUFCMINSTRUCTION(17),
	GlitchData    => APUFCMINSTRUCTION17_GlitchData,
	OutSignalName => "APUFCMINSTRUCTION(17)",
	OutTemp       => APUFCMINSTRUCTION_OUT(17),
	Paths         => (0 => (CPMFCMCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => APUFCMINSTRUCTION(18),
	GlitchData    => APUFCMINSTRUCTION18_GlitchData,
	OutSignalName => "APUFCMINSTRUCTION(18)",
	OutTemp       => APUFCMINSTRUCTION_OUT(18),
	Paths         => (0 => (CPMFCMCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => APUFCMINSTRUCTION(19),
	GlitchData    => APUFCMINSTRUCTION19_GlitchData,
	OutSignalName => "APUFCMINSTRUCTION(19)",
	OutTemp       => APUFCMINSTRUCTION_OUT(19),
	Paths         => (0 => (CPMFCMCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => APUFCMINSTRUCTION(20),
	GlitchData    => APUFCMINSTRUCTION20_GlitchData,
	OutSignalName => "APUFCMINSTRUCTION(20)",
	OutTemp       => APUFCMINSTRUCTION_OUT(20),
	Paths         => (0 => (CPMFCMCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => APUFCMINSTRUCTION(21),
	GlitchData    => APUFCMINSTRUCTION21_GlitchData,
	OutSignalName => "APUFCMINSTRUCTION(21)",
	OutTemp       => APUFCMINSTRUCTION_OUT(21),
	Paths         => (0 => (CPMFCMCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => APUFCMINSTRUCTION(22),
	GlitchData    => APUFCMINSTRUCTION22_GlitchData,
	OutSignalName => "APUFCMINSTRUCTION(22)",
	OutTemp       => APUFCMINSTRUCTION_OUT(22),
	Paths         => (0 => (CPMFCMCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => APUFCMINSTRUCTION(23),
	GlitchData    => APUFCMINSTRUCTION23_GlitchData,
	OutSignalName => "APUFCMINSTRUCTION(23)",
	OutTemp       => APUFCMINSTRUCTION_OUT(23),
	Paths         => (0 => (CPMFCMCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => APUFCMINSTRUCTION(24),
	GlitchData    => APUFCMINSTRUCTION24_GlitchData,
	OutSignalName => "APUFCMINSTRUCTION(24)",
	OutTemp       => APUFCMINSTRUCTION_OUT(24),
	Paths         => (0 => (CPMFCMCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => APUFCMINSTRUCTION(25),
	GlitchData    => APUFCMINSTRUCTION25_GlitchData,
	OutSignalName => "APUFCMINSTRUCTION(25)",
	OutTemp       => APUFCMINSTRUCTION_OUT(25),
	Paths         => (0 => (CPMFCMCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => APUFCMINSTRUCTION(26),
	GlitchData    => APUFCMINSTRUCTION26_GlitchData,
	OutSignalName => "APUFCMINSTRUCTION(26)",
	OutTemp       => APUFCMINSTRUCTION_OUT(26),
	Paths         => (0 => (CPMFCMCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => APUFCMINSTRUCTION(27),
	GlitchData    => APUFCMINSTRUCTION27_GlitchData,
	OutSignalName => "APUFCMINSTRUCTION(27)",
	OutTemp       => APUFCMINSTRUCTION_OUT(27),
	Paths         => (0 => (CPMFCMCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => APUFCMINSTRUCTION(28),
	GlitchData    => APUFCMINSTRUCTION28_GlitchData,
	OutSignalName => "APUFCMINSTRUCTION(28)",
	OutTemp       => APUFCMINSTRUCTION_OUT(28),
	Paths         => (0 => (CPMFCMCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => APUFCMINSTRUCTION(29),
	GlitchData    => APUFCMINSTRUCTION29_GlitchData,
	OutSignalName => "APUFCMINSTRUCTION(29)",
	OutTemp       => APUFCMINSTRUCTION_OUT(29),
	Paths         => (0 => (CPMFCMCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => APUFCMINSTRUCTION(30),
	GlitchData    => APUFCMINSTRUCTION30_GlitchData,
	OutSignalName => "APUFCMINSTRUCTION(30)",
	OutTemp       => APUFCMINSTRUCTION_OUT(30),
	Paths         => (0 => (CPMFCMCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => APUFCMINSTRUCTION(31),
	GlitchData    => APUFCMINSTRUCTION31_GlitchData,
	OutSignalName => "APUFCMINSTRUCTION(31)",
	OutTemp       => APUFCMINSTRUCTION_OUT(31),
	Paths         => (0 => (CPMFCMCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => APUFCMINSTRVALID,
	GlitchData    => APUFCMINSTRVALID_GlitchData,
	OutSignalName => "APUFCMINSTRVALID",
	OutTemp       => APUFCMINSTRVALID_OUT,
	Paths         => (0 => (CPMFCMCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => APUFCMLOADBYTEADDR(0),
	GlitchData    => APUFCMLOADBYTEADDR0_GlitchData,
	OutSignalName => "APUFCMLOADBYTEADDR(0)",
	OutTemp       => APUFCMLOADBYTEADDR_OUT(0),
	Paths         => (0 => (CPMFCMCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => APUFCMLOADBYTEADDR(1),
	GlitchData    => APUFCMLOADBYTEADDR1_GlitchData,
	OutSignalName => "APUFCMLOADBYTEADDR(1)",
	OutTemp       => APUFCMLOADBYTEADDR_OUT(1),
	Paths         => (0 => (CPMFCMCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => APUFCMLOADBYTEADDR(2),
	GlitchData    => APUFCMLOADBYTEADDR2_GlitchData,
	OutSignalName => "APUFCMLOADBYTEADDR(2)",
	OutTemp       => APUFCMLOADBYTEADDR_OUT(2),
	Paths         => (0 => (CPMFCMCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => APUFCMLOADBYTEADDR(3),
	GlitchData    => APUFCMLOADBYTEADDR3_GlitchData,
	OutSignalName => "APUFCMLOADBYTEADDR(3)",
	OutTemp       => APUFCMLOADBYTEADDR_OUT(3),
	Paths         => (0 => (CPMFCMCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => APUFCMLOADDATA(0),
	GlitchData    => APUFCMLOADDATA0_GlitchData,
	OutSignalName => "APUFCMLOADDATA(0)",
	OutTemp       => APUFCMLOADDATA_OUT(0),
	Paths         => (0 => (CPMFCMCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => APUFCMLOADDATA(1),
	GlitchData    => APUFCMLOADDATA1_GlitchData,
	OutSignalName => "APUFCMLOADDATA(1)",
	OutTemp       => APUFCMLOADDATA_OUT(1),
	Paths         => (0 => (CPMFCMCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => APUFCMLOADDATA(2),
	GlitchData    => APUFCMLOADDATA2_GlitchData,
	OutSignalName => "APUFCMLOADDATA(2)",
	OutTemp       => APUFCMLOADDATA_OUT(2),
	Paths         => (0 => (CPMFCMCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => APUFCMLOADDATA(3),
	GlitchData    => APUFCMLOADDATA3_GlitchData,
	OutSignalName => "APUFCMLOADDATA(3)",
	OutTemp       => APUFCMLOADDATA_OUT(3),
	Paths         => (0 => (CPMFCMCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => APUFCMLOADDATA(4),
	GlitchData    => APUFCMLOADDATA4_GlitchData,
	OutSignalName => "APUFCMLOADDATA(4)",
	OutTemp       => APUFCMLOADDATA_OUT(4),
	Paths         => (0 => (CPMFCMCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => APUFCMLOADDATA(5),
	GlitchData    => APUFCMLOADDATA5_GlitchData,
	OutSignalName => "APUFCMLOADDATA(5)",
	OutTemp       => APUFCMLOADDATA_OUT(5),
	Paths         => (0 => (CPMFCMCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => APUFCMLOADDATA(6),
	GlitchData    => APUFCMLOADDATA6_GlitchData,
	OutSignalName => "APUFCMLOADDATA(6)",
	OutTemp       => APUFCMLOADDATA_OUT(6),
	Paths         => (0 => (CPMFCMCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => APUFCMLOADDATA(7),
	GlitchData    => APUFCMLOADDATA7_GlitchData,
	OutSignalName => "APUFCMLOADDATA(7)",
	OutTemp       => APUFCMLOADDATA_OUT(7),
	Paths         => (0 => (CPMFCMCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => APUFCMLOADDATA(8),
	GlitchData    => APUFCMLOADDATA8_GlitchData,
	OutSignalName => "APUFCMLOADDATA(8)",
	OutTemp       => APUFCMLOADDATA_OUT(8),
	Paths         => (0 => (CPMFCMCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => APUFCMLOADDATA(9),
	GlitchData    => APUFCMLOADDATA9_GlitchData,
	OutSignalName => "APUFCMLOADDATA(9)",
	OutTemp       => APUFCMLOADDATA_OUT(9),
	Paths         => (0 => (CPMFCMCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => APUFCMLOADDATA(10),
	GlitchData    => APUFCMLOADDATA10_GlitchData,
	OutSignalName => "APUFCMLOADDATA(10)",
	OutTemp       => APUFCMLOADDATA_OUT(10),
	Paths         => (0 => (CPMFCMCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => APUFCMLOADDATA(11),
	GlitchData    => APUFCMLOADDATA11_GlitchData,
	OutSignalName => "APUFCMLOADDATA(11)",
	OutTemp       => APUFCMLOADDATA_OUT(11),
	Paths         => (0 => (CPMFCMCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => APUFCMLOADDATA(12),
	GlitchData    => APUFCMLOADDATA12_GlitchData,
	OutSignalName => "APUFCMLOADDATA(12)",
	OutTemp       => APUFCMLOADDATA_OUT(12),
	Paths         => (0 => (CPMFCMCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => APUFCMLOADDATA(13),
	GlitchData    => APUFCMLOADDATA13_GlitchData,
	OutSignalName => "APUFCMLOADDATA(13)",
	OutTemp       => APUFCMLOADDATA_OUT(13),
	Paths         => (0 => (CPMFCMCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => APUFCMLOADDATA(14),
	GlitchData    => APUFCMLOADDATA14_GlitchData,
	OutSignalName => "APUFCMLOADDATA(14)",
	OutTemp       => APUFCMLOADDATA_OUT(14),
	Paths         => (0 => (CPMFCMCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => APUFCMLOADDATA(15),
	GlitchData    => APUFCMLOADDATA15_GlitchData,
	OutSignalName => "APUFCMLOADDATA(15)",
	OutTemp       => APUFCMLOADDATA_OUT(15),
	Paths         => (0 => (CPMFCMCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => APUFCMLOADDATA(16),
	GlitchData    => APUFCMLOADDATA16_GlitchData,
	OutSignalName => "APUFCMLOADDATA(16)",
	OutTemp       => APUFCMLOADDATA_OUT(16),
	Paths         => (0 => (CPMFCMCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => APUFCMLOADDATA(17),
	GlitchData    => APUFCMLOADDATA17_GlitchData,
	OutSignalName => "APUFCMLOADDATA(17)",
	OutTemp       => APUFCMLOADDATA_OUT(17),
	Paths         => (0 => (CPMFCMCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => APUFCMLOADDATA(18),
	GlitchData    => APUFCMLOADDATA18_GlitchData,
	OutSignalName => "APUFCMLOADDATA(18)",
	OutTemp       => APUFCMLOADDATA_OUT(18),
	Paths         => (0 => (CPMFCMCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => APUFCMLOADDATA(19),
	GlitchData    => APUFCMLOADDATA19_GlitchData,
	OutSignalName => "APUFCMLOADDATA(19)",
	OutTemp       => APUFCMLOADDATA_OUT(19),
	Paths         => (0 => (CPMFCMCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => APUFCMLOADDATA(20),
	GlitchData    => APUFCMLOADDATA20_GlitchData,
	OutSignalName => "APUFCMLOADDATA(20)",
	OutTemp       => APUFCMLOADDATA_OUT(20),
	Paths         => (0 => (CPMFCMCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => APUFCMLOADDATA(21),
	GlitchData    => APUFCMLOADDATA21_GlitchData,
	OutSignalName => "APUFCMLOADDATA(21)",
	OutTemp       => APUFCMLOADDATA_OUT(21),
	Paths         => (0 => (CPMFCMCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => APUFCMLOADDATA(22),
	GlitchData    => APUFCMLOADDATA22_GlitchData,
	OutSignalName => "APUFCMLOADDATA(22)",
	OutTemp       => APUFCMLOADDATA_OUT(22),
	Paths         => (0 => (CPMFCMCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => APUFCMLOADDATA(23),
	GlitchData    => APUFCMLOADDATA23_GlitchData,
	OutSignalName => "APUFCMLOADDATA(23)",
	OutTemp       => APUFCMLOADDATA_OUT(23),
	Paths         => (0 => (CPMFCMCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => APUFCMLOADDATA(24),
	GlitchData    => APUFCMLOADDATA24_GlitchData,
	OutSignalName => "APUFCMLOADDATA(24)",
	OutTemp       => APUFCMLOADDATA_OUT(24),
	Paths         => (0 => (CPMFCMCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => APUFCMLOADDATA(25),
	GlitchData    => APUFCMLOADDATA25_GlitchData,
	OutSignalName => "APUFCMLOADDATA(25)",
	OutTemp       => APUFCMLOADDATA_OUT(25),
	Paths         => (0 => (CPMFCMCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => APUFCMLOADDATA(26),
	GlitchData    => APUFCMLOADDATA26_GlitchData,
	OutSignalName => "APUFCMLOADDATA(26)",
	OutTemp       => APUFCMLOADDATA_OUT(26),
	Paths         => (0 => (CPMFCMCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => APUFCMLOADDATA(27),
	GlitchData    => APUFCMLOADDATA27_GlitchData,
	OutSignalName => "APUFCMLOADDATA(27)",
	OutTemp       => APUFCMLOADDATA_OUT(27),
	Paths         => (0 => (CPMFCMCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => APUFCMLOADDATA(28),
	GlitchData    => APUFCMLOADDATA28_GlitchData,
	OutSignalName => "APUFCMLOADDATA(28)",
	OutTemp       => APUFCMLOADDATA_OUT(28),
	Paths         => (0 => (CPMFCMCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => APUFCMLOADDATA(29),
	GlitchData    => APUFCMLOADDATA29_GlitchData,
	OutSignalName => "APUFCMLOADDATA(29)",
	OutTemp       => APUFCMLOADDATA_OUT(29),
	Paths         => (0 => (CPMFCMCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => APUFCMLOADDATA(30),
	GlitchData    => APUFCMLOADDATA30_GlitchData,
	OutSignalName => "APUFCMLOADDATA(30)",
	OutTemp       => APUFCMLOADDATA_OUT(30),
	Paths         => (0 => (CPMFCMCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => APUFCMLOADDATA(31),
	GlitchData    => APUFCMLOADDATA31_GlitchData,
	OutSignalName => "APUFCMLOADDATA(31)",
	OutTemp       => APUFCMLOADDATA_OUT(31),
	Paths         => (0 => (CPMFCMCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => APUFCMLOADDATA(32),
	GlitchData    => APUFCMLOADDATA32_GlitchData,
	OutSignalName => "APUFCMLOADDATA(32)",
	OutTemp       => APUFCMLOADDATA_OUT(32),
	Paths         => (0 => (CPMFCMCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => APUFCMLOADDATA(33),
	GlitchData    => APUFCMLOADDATA33_GlitchData,
	OutSignalName => "APUFCMLOADDATA(33)",
	OutTemp       => APUFCMLOADDATA_OUT(33),
	Paths         => (0 => (CPMFCMCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => APUFCMLOADDATA(34),
	GlitchData    => APUFCMLOADDATA34_GlitchData,
	OutSignalName => "APUFCMLOADDATA(34)",
	OutTemp       => APUFCMLOADDATA_OUT(34),
	Paths         => (0 => (CPMFCMCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => APUFCMLOADDATA(35),
	GlitchData    => APUFCMLOADDATA35_GlitchData,
	OutSignalName => "APUFCMLOADDATA(35)",
	OutTemp       => APUFCMLOADDATA_OUT(35),
	Paths         => (0 => (CPMFCMCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => APUFCMLOADDATA(36),
	GlitchData    => APUFCMLOADDATA36_GlitchData,
	OutSignalName => "APUFCMLOADDATA(36)",
	OutTemp       => APUFCMLOADDATA_OUT(36),
	Paths         => (0 => (CPMFCMCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => APUFCMLOADDATA(37),
	GlitchData    => APUFCMLOADDATA37_GlitchData,
	OutSignalName => "APUFCMLOADDATA(37)",
	OutTemp       => APUFCMLOADDATA_OUT(37),
	Paths         => (0 => (CPMFCMCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => APUFCMLOADDATA(38),
	GlitchData    => APUFCMLOADDATA38_GlitchData,
	OutSignalName => "APUFCMLOADDATA(38)",
	OutTemp       => APUFCMLOADDATA_OUT(38),
	Paths         => (0 => (CPMFCMCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => APUFCMLOADDATA(39),
	GlitchData    => APUFCMLOADDATA39_GlitchData,
	OutSignalName => "APUFCMLOADDATA(39)",
	OutTemp       => APUFCMLOADDATA_OUT(39),
	Paths         => (0 => (CPMFCMCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => APUFCMLOADDATA(40),
	GlitchData    => APUFCMLOADDATA40_GlitchData,
	OutSignalName => "APUFCMLOADDATA(40)",
	OutTemp       => APUFCMLOADDATA_OUT(40),
	Paths         => (0 => (CPMFCMCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => APUFCMLOADDATA(41),
	GlitchData    => APUFCMLOADDATA41_GlitchData,
	OutSignalName => "APUFCMLOADDATA(41)",
	OutTemp       => APUFCMLOADDATA_OUT(41),
	Paths         => (0 => (CPMFCMCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => APUFCMLOADDATA(42),
	GlitchData    => APUFCMLOADDATA42_GlitchData,
	OutSignalName => "APUFCMLOADDATA(42)",
	OutTemp       => APUFCMLOADDATA_OUT(42),
	Paths         => (0 => (CPMFCMCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => APUFCMLOADDATA(43),
	GlitchData    => APUFCMLOADDATA43_GlitchData,
	OutSignalName => "APUFCMLOADDATA(43)",
	OutTemp       => APUFCMLOADDATA_OUT(43),
	Paths         => (0 => (CPMFCMCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => APUFCMLOADDATA(44),
	GlitchData    => APUFCMLOADDATA44_GlitchData,
	OutSignalName => "APUFCMLOADDATA(44)",
	OutTemp       => APUFCMLOADDATA_OUT(44),
	Paths         => (0 => (CPMFCMCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => APUFCMLOADDATA(45),
	GlitchData    => APUFCMLOADDATA45_GlitchData,
	OutSignalName => "APUFCMLOADDATA(45)",
	OutTemp       => APUFCMLOADDATA_OUT(45),
	Paths         => (0 => (CPMFCMCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => APUFCMLOADDATA(46),
	GlitchData    => APUFCMLOADDATA46_GlitchData,
	OutSignalName => "APUFCMLOADDATA(46)",
	OutTemp       => APUFCMLOADDATA_OUT(46),
	Paths         => (0 => (CPMFCMCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => APUFCMLOADDATA(47),
	GlitchData    => APUFCMLOADDATA47_GlitchData,
	OutSignalName => "APUFCMLOADDATA(47)",
	OutTemp       => APUFCMLOADDATA_OUT(47),
	Paths         => (0 => (CPMFCMCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => APUFCMLOADDATA(48),
	GlitchData    => APUFCMLOADDATA48_GlitchData,
	OutSignalName => "APUFCMLOADDATA(48)",
	OutTemp       => APUFCMLOADDATA_OUT(48),
	Paths         => (0 => (CPMFCMCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => APUFCMLOADDATA(49),
	GlitchData    => APUFCMLOADDATA49_GlitchData,
	OutSignalName => "APUFCMLOADDATA(49)",
	OutTemp       => APUFCMLOADDATA_OUT(49),
	Paths         => (0 => (CPMFCMCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => APUFCMLOADDATA(50),
	GlitchData    => APUFCMLOADDATA50_GlitchData,
	OutSignalName => "APUFCMLOADDATA(50)",
	OutTemp       => APUFCMLOADDATA_OUT(50),
	Paths         => (0 => (CPMFCMCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => APUFCMLOADDATA(51),
	GlitchData    => APUFCMLOADDATA51_GlitchData,
	OutSignalName => "APUFCMLOADDATA(51)",
	OutTemp       => APUFCMLOADDATA_OUT(51),
	Paths         => (0 => (CPMFCMCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => APUFCMLOADDATA(52),
	GlitchData    => APUFCMLOADDATA52_GlitchData,
	OutSignalName => "APUFCMLOADDATA(52)",
	OutTemp       => APUFCMLOADDATA_OUT(52),
	Paths         => (0 => (CPMFCMCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => APUFCMLOADDATA(53),
	GlitchData    => APUFCMLOADDATA53_GlitchData,
	OutSignalName => "APUFCMLOADDATA(53)",
	OutTemp       => APUFCMLOADDATA_OUT(53),
	Paths         => (0 => (CPMFCMCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => APUFCMLOADDATA(54),
	GlitchData    => APUFCMLOADDATA54_GlitchData,
	OutSignalName => "APUFCMLOADDATA(54)",
	OutTemp       => APUFCMLOADDATA_OUT(54),
	Paths         => (0 => (CPMFCMCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => APUFCMLOADDATA(55),
	GlitchData    => APUFCMLOADDATA55_GlitchData,
	OutSignalName => "APUFCMLOADDATA(55)",
	OutTemp       => APUFCMLOADDATA_OUT(55),
	Paths         => (0 => (CPMFCMCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => APUFCMLOADDATA(56),
	GlitchData    => APUFCMLOADDATA56_GlitchData,
	OutSignalName => "APUFCMLOADDATA(56)",
	OutTemp       => APUFCMLOADDATA_OUT(56),
	Paths         => (0 => (CPMFCMCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => APUFCMLOADDATA(57),
	GlitchData    => APUFCMLOADDATA57_GlitchData,
	OutSignalName => "APUFCMLOADDATA(57)",
	OutTemp       => APUFCMLOADDATA_OUT(57),
	Paths         => (0 => (CPMFCMCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => APUFCMLOADDATA(58),
	GlitchData    => APUFCMLOADDATA58_GlitchData,
	OutSignalName => "APUFCMLOADDATA(58)",
	OutTemp       => APUFCMLOADDATA_OUT(58),
	Paths         => (0 => (CPMFCMCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => APUFCMLOADDATA(59),
	GlitchData    => APUFCMLOADDATA59_GlitchData,
	OutSignalName => "APUFCMLOADDATA(59)",
	OutTemp       => APUFCMLOADDATA_OUT(59),
	Paths         => (0 => (CPMFCMCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => APUFCMLOADDATA(60),
	GlitchData    => APUFCMLOADDATA60_GlitchData,
	OutSignalName => "APUFCMLOADDATA(60)",
	OutTemp       => APUFCMLOADDATA_OUT(60),
	Paths         => (0 => (CPMFCMCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => APUFCMLOADDATA(61),
	GlitchData    => APUFCMLOADDATA61_GlitchData,
	OutSignalName => "APUFCMLOADDATA(61)",
	OutTemp       => APUFCMLOADDATA_OUT(61),
	Paths         => (0 => (CPMFCMCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => APUFCMLOADDATA(62),
	GlitchData    => APUFCMLOADDATA62_GlitchData,
	OutSignalName => "APUFCMLOADDATA(62)",
	OutTemp       => APUFCMLOADDATA_OUT(62),
	Paths         => (0 => (CPMFCMCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => APUFCMLOADDATA(63),
	GlitchData    => APUFCMLOADDATA63_GlitchData,
	OutSignalName => "APUFCMLOADDATA(63)",
	OutTemp       => APUFCMLOADDATA_OUT(63),
	Paths         => (0 => (CPMFCMCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => APUFCMLOADDATA(64),
	GlitchData    => APUFCMLOADDATA64_GlitchData,
	OutSignalName => "APUFCMLOADDATA(64)",
	OutTemp       => APUFCMLOADDATA_OUT(64),
	Paths         => (0 => (CPMFCMCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => APUFCMLOADDATA(65),
	GlitchData    => APUFCMLOADDATA65_GlitchData,
	OutSignalName => "APUFCMLOADDATA(65)",
	OutTemp       => APUFCMLOADDATA_OUT(65),
	Paths         => (0 => (CPMFCMCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => APUFCMLOADDATA(66),
	GlitchData    => APUFCMLOADDATA66_GlitchData,
	OutSignalName => "APUFCMLOADDATA(66)",
	OutTemp       => APUFCMLOADDATA_OUT(66),
	Paths         => (0 => (CPMFCMCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => APUFCMLOADDATA(67),
	GlitchData    => APUFCMLOADDATA67_GlitchData,
	OutSignalName => "APUFCMLOADDATA(67)",
	OutTemp       => APUFCMLOADDATA_OUT(67),
	Paths         => (0 => (CPMFCMCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => APUFCMLOADDATA(68),
	GlitchData    => APUFCMLOADDATA68_GlitchData,
	OutSignalName => "APUFCMLOADDATA(68)",
	OutTemp       => APUFCMLOADDATA_OUT(68),
	Paths         => (0 => (CPMFCMCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => APUFCMLOADDATA(69),
	GlitchData    => APUFCMLOADDATA69_GlitchData,
	OutSignalName => "APUFCMLOADDATA(69)",
	OutTemp       => APUFCMLOADDATA_OUT(69),
	Paths         => (0 => (CPMFCMCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => APUFCMLOADDATA(70),
	GlitchData    => APUFCMLOADDATA70_GlitchData,
	OutSignalName => "APUFCMLOADDATA(70)",
	OutTemp       => APUFCMLOADDATA_OUT(70),
	Paths         => (0 => (CPMFCMCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => APUFCMLOADDATA(71),
	GlitchData    => APUFCMLOADDATA71_GlitchData,
	OutSignalName => "APUFCMLOADDATA(71)",
	OutTemp       => APUFCMLOADDATA_OUT(71),
	Paths         => (0 => (CPMFCMCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => APUFCMLOADDATA(72),
	GlitchData    => APUFCMLOADDATA72_GlitchData,
	OutSignalName => "APUFCMLOADDATA(72)",
	OutTemp       => APUFCMLOADDATA_OUT(72),
	Paths         => (0 => (CPMFCMCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => APUFCMLOADDATA(73),
	GlitchData    => APUFCMLOADDATA73_GlitchData,
	OutSignalName => "APUFCMLOADDATA(73)",
	OutTemp       => APUFCMLOADDATA_OUT(73),
	Paths         => (0 => (CPMFCMCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => APUFCMLOADDATA(74),
	GlitchData    => APUFCMLOADDATA74_GlitchData,
	OutSignalName => "APUFCMLOADDATA(74)",
	OutTemp       => APUFCMLOADDATA_OUT(74),
	Paths         => (0 => (CPMFCMCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => APUFCMLOADDATA(75),
	GlitchData    => APUFCMLOADDATA75_GlitchData,
	OutSignalName => "APUFCMLOADDATA(75)",
	OutTemp       => APUFCMLOADDATA_OUT(75),
	Paths         => (0 => (CPMFCMCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => APUFCMLOADDATA(76),
	GlitchData    => APUFCMLOADDATA76_GlitchData,
	OutSignalName => "APUFCMLOADDATA(76)",
	OutTemp       => APUFCMLOADDATA_OUT(76),
	Paths         => (0 => (CPMFCMCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => APUFCMLOADDATA(77),
	GlitchData    => APUFCMLOADDATA77_GlitchData,
	OutSignalName => "APUFCMLOADDATA(77)",
	OutTemp       => APUFCMLOADDATA_OUT(77),
	Paths         => (0 => (CPMFCMCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => APUFCMLOADDATA(78),
	GlitchData    => APUFCMLOADDATA78_GlitchData,
	OutSignalName => "APUFCMLOADDATA(78)",
	OutTemp       => APUFCMLOADDATA_OUT(78),
	Paths         => (0 => (CPMFCMCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => APUFCMLOADDATA(79),
	GlitchData    => APUFCMLOADDATA79_GlitchData,
	OutSignalName => "APUFCMLOADDATA(79)",
	OutTemp       => APUFCMLOADDATA_OUT(79),
	Paths         => (0 => (CPMFCMCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => APUFCMLOADDATA(80),
	GlitchData    => APUFCMLOADDATA80_GlitchData,
	OutSignalName => "APUFCMLOADDATA(80)",
	OutTemp       => APUFCMLOADDATA_OUT(80),
	Paths         => (0 => (CPMFCMCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => APUFCMLOADDATA(81),
	GlitchData    => APUFCMLOADDATA81_GlitchData,
	OutSignalName => "APUFCMLOADDATA(81)",
	OutTemp       => APUFCMLOADDATA_OUT(81),
	Paths         => (0 => (CPMFCMCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => APUFCMLOADDATA(82),
	GlitchData    => APUFCMLOADDATA82_GlitchData,
	OutSignalName => "APUFCMLOADDATA(82)",
	OutTemp       => APUFCMLOADDATA_OUT(82),
	Paths         => (0 => (CPMFCMCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => APUFCMLOADDATA(83),
	GlitchData    => APUFCMLOADDATA83_GlitchData,
	OutSignalName => "APUFCMLOADDATA(83)",
	OutTemp       => APUFCMLOADDATA_OUT(83),
	Paths         => (0 => (CPMFCMCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => APUFCMLOADDATA(84),
	GlitchData    => APUFCMLOADDATA84_GlitchData,
	OutSignalName => "APUFCMLOADDATA(84)",
	OutTemp       => APUFCMLOADDATA_OUT(84),
	Paths         => (0 => (CPMFCMCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => APUFCMLOADDATA(85),
	GlitchData    => APUFCMLOADDATA85_GlitchData,
	OutSignalName => "APUFCMLOADDATA(85)",
	OutTemp       => APUFCMLOADDATA_OUT(85),
	Paths         => (0 => (CPMFCMCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => APUFCMLOADDATA(86),
	GlitchData    => APUFCMLOADDATA86_GlitchData,
	OutSignalName => "APUFCMLOADDATA(86)",
	OutTemp       => APUFCMLOADDATA_OUT(86),
	Paths         => (0 => (CPMFCMCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => APUFCMLOADDATA(87),
	GlitchData    => APUFCMLOADDATA87_GlitchData,
	OutSignalName => "APUFCMLOADDATA(87)",
	OutTemp       => APUFCMLOADDATA_OUT(87),
	Paths         => (0 => (CPMFCMCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => APUFCMLOADDATA(88),
	GlitchData    => APUFCMLOADDATA88_GlitchData,
	OutSignalName => "APUFCMLOADDATA(88)",
	OutTemp       => APUFCMLOADDATA_OUT(88),
	Paths         => (0 => (CPMFCMCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => APUFCMLOADDATA(89),
	GlitchData    => APUFCMLOADDATA89_GlitchData,
	OutSignalName => "APUFCMLOADDATA(89)",
	OutTemp       => APUFCMLOADDATA_OUT(89),
	Paths         => (0 => (CPMFCMCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => APUFCMLOADDATA(90),
	GlitchData    => APUFCMLOADDATA90_GlitchData,
	OutSignalName => "APUFCMLOADDATA(90)",
	OutTemp       => APUFCMLOADDATA_OUT(90),
	Paths         => (0 => (CPMFCMCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => APUFCMLOADDATA(91),
	GlitchData    => APUFCMLOADDATA91_GlitchData,
	OutSignalName => "APUFCMLOADDATA(91)",
	OutTemp       => APUFCMLOADDATA_OUT(91),
	Paths         => (0 => (CPMFCMCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => APUFCMLOADDATA(92),
	GlitchData    => APUFCMLOADDATA92_GlitchData,
	OutSignalName => "APUFCMLOADDATA(92)",
	OutTemp       => APUFCMLOADDATA_OUT(92),
	Paths         => (0 => (CPMFCMCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => APUFCMLOADDATA(93),
	GlitchData    => APUFCMLOADDATA93_GlitchData,
	OutSignalName => "APUFCMLOADDATA(93)",
	OutTemp       => APUFCMLOADDATA_OUT(93),
	Paths         => (0 => (CPMFCMCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => APUFCMLOADDATA(94),
	GlitchData    => APUFCMLOADDATA94_GlitchData,
	OutSignalName => "APUFCMLOADDATA(94)",
	OutTemp       => APUFCMLOADDATA_OUT(94),
	Paths         => (0 => (CPMFCMCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => APUFCMLOADDATA(95),
	GlitchData    => APUFCMLOADDATA95_GlitchData,
	OutSignalName => "APUFCMLOADDATA(95)",
	OutTemp       => APUFCMLOADDATA_OUT(95),
	Paths         => (0 => (CPMFCMCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => APUFCMLOADDATA(96),
	GlitchData    => APUFCMLOADDATA96_GlitchData,
	OutSignalName => "APUFCMLOADDATA(96)",
	OutTemp       => APUFCMLOADDATA_OUT(96),
	Paths         => (0 => (CPMFCMCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => APUFCMLOADDATA(97),
	GlitchData    => APUFCMLOADDATA97_GlitchData,
	OutSignalName => "APUFCMLOADDATA(97)",
	OutTemp       => APUFCMLOADDATA_OUT(97),
	Paths         => (0 => (CPMFCMCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => APUFCMLOADDATA(98),
	GlitchData    => APUFCMLOADDATA98_GlitchData,
	OutSignalName => "APUFCMLOADDATA(98)",
	OutTemp       => APUFCMLOADDATA_OUT(98),
	Paths         => (0 => (CPMFCMCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => APUFCMLOADDATA(99),
	GlitchData    => APUFCMLOADDATA99_GlitchData,
	OutSignalName => "APUFCMLOADDATA(99)",
	OutTemp       => APUFCMLOADDATA_OUT(99),
	Paths         => (0 => (CPMFCMCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => APUFCMLOADDATA(100),
	GlitchData    => APUFCMLOADDATA100_GlitchData,
	OutSignalName => "APUFCMLOADDATA(100)",
	OutTemp       => APUFCMLOADDATA_OUT(100),
	Paths         => (0 => (CPMFCMCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => APUFCMLOADDATA(101),
	GlitchData    => APUFCMLOADDATA101_GlitchData,
	OutSignalName => "APUFCMLOADDATA(101)",
	OutTemp       => APUFCMLOADDATA_OUT(101),
	Paths         => (0 => (CPMFCMCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => APUFCMLOADDATA(102),
	GlitchData    => APUFCMLOADDATA102_GlitchData,
	OutSignalName => "APUFCMLOADDATA(102)",
	OutTemp       => APUFCMLOADDATA_OUT(102),
	Paths         => (0 => (CPMFCMCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => APUFCMLOADDATA(103),
	GlitchData    => APUFCMLOADDATA103_GlitchData,
	OutSignalName => "APUFCMLOADDATA(103)",
	OutTemp       => APUFCMLOADDATA_OUT(103),
	Paths         => (0 => (CPMFCMCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => APUFCMLOADDATA(104),
	GlitchData    => APUFCMLOADDATA104_GlitchData,
	OutSignalName => "APUFCMLOADDATA(104)",
	OutTemp       => APUFCMLOADDATA_OUT(104),
	Paths         => (0 => (CPMFCMCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => APUFCMLOADDATA(105),
	GlitchData    => APUFCMLOADDATA105_GlitchData,
	OutSignalName => "APUFCMLOADDATA(105)",
	OutTemp       => APUFCMLOADDATA_OUT(105),
	Paths         => (0 => (CPMFCMCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => APUFCMLOADDATA(106),
	GlitchData    => APUFCMLOADDATA106_GlitchData,
	OutSignalName => "APUFCMLOADDATA(106)",
	OutTemp       => APUFCMLOADDATA_OUT(106),
	Paths         => (0 => (CPMFCMCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => APUFCMLOADDATA(107),
	GlitchData    => APUFCMLOADDATA107_GlitchData,
	OutSignalName => "APUFCMLOADDATA(107)",
	OutTemp       => APUFCMLOADDATA_OUT(107),
	Paths         => (0 => (CPMFCMCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => APUFCMLOADDATA(108),
	GlitchData    => APUFCMLOADDATA108_GlitchData,
	OutSignalName => "APUFCMLOADDATA(108)",
	OutTemp       => APUFCMLOADDATA_OUT(108),
	Paths         => (0 => (CPMFCMCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => APUFCMLOADDATA(109),
	GlitchData    => APUFCMLOADDATA109_GlitchData,
	OutSignalName => "APUFCMLOADDATA(109)",
	OutTemp       => APUFCMLOADDATA_OUT(109),
	Paths         => (0 => (CPMFCMCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => APUFCMLOADDATA(110),
	GlitchData    => APUFCMLOADDATA110_GlitchData,
	OutSignalName => "APUFCMLOADDATA(110)",
	OutTemp       => APUFCMLOADDATA_OUT(110),
	Paths         => (0 => (CPMFCMCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => APUFCMLOADDATA(111),
	GlitchData    => APUFCMLOADDATA111_GlitchData,
	OutSignalName => "APUFCMLOADDATA(111)",
	OutTemp       => APUFCMLOADDATA_OUT(111),
	Paths         => (0 => (CPMFCMCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => APUFCMLOADDATA(112),
	GlitchData    => APUFCMLOADDATA112_GlitchData,
	OutSignalName => "APUFCMLOADDATA(112)",
	OutTemp       => APUFCMLOADDATA_OUT(112),
	Paths         => (0 => (CPMFCMCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => APUFCMLOADDATA(113),
	GlitchData    => APUFCMLOADDATA113_GlitchData,
	OutSignalName => "APUFCMLOADDATA(113)",
	OutTemp       => APUFCMLOADDATA_OUT(113),
	Paths         => (0 => (CPMFCMCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => APUFCMLOADDATA(114),
	GlitchData    => APUFCMLOADDATA114_GlitchData,
	OutSignalName => "APUFCMLOADDATA(114)",
	OutTemp       => APUFCMLOADDATA_OUT(114),
	Paths         => (0 => (CPMFCMCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => APUFCMLOADDATA(115),
	GlitchData    => APUFCMLOADDATA115_GlitchData,
	OutSignalName => "APUFCMLOADDATA(115)",
	OutTemp       => APUFCMLOADDATA_OUT(115),
	Paths         => (0 => (CPMFCMCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => APUFCMLOADDATA(116),
	GlitchData    => APUFCMLOADDATA116_GlitchData,
	OutSignalName => "APUFCMLOADDATA(116)",
	OutTemp       => APUFCMLOADDATA_OUT(116),
	Paths         => (0 => (CPMFCMCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => APUFCMLOADDATA(117),
	GlitchData    => APUFCMLOADDATA117_GlitchData,
	OutSignalName => "APUFCMLOADDATA(117)",
	OutTemp       => APUFCMLOADDATA_OUT(117),
	Paths         => (0 => (CPMFCMCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => APUFCMLOADDATA(118),
	GlitchData    => APUFCMLOADDATA118_GlitchData,
	OutSignalName => "APUFCMLOADDATA(118)",
	OutTemp       => APUFCMLOADDATA_OUT(118),
	Paths         => (0 => (CPMFCMCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => APUFCMLOADDATA(119),
	GlitchData    => APUFCMLOADDATA119_GlitchData,
	OutSignalName => "APUFCMLOADDATA(119)",
	OutTemp       => APUFCMLOADDATA_OUT(119),
	Paths         => (0 => (CPMFCMCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => APUFCMLOADDATA(120),
	GlitchData    => APUFCMLOADDATA120_GlitchData,
	OutSignalName => "APUFCMLOADDATA(120)",
	OutTemp       => APUFCMLOADDATA_OUT(120),
	Paths         => (0 => (CPMFCMCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => APUFCMLOADDATA(121),
	GlitchData    => APUFCMLOADDATA121_GlitchData,
	OutSignalName => "APUFCMLOADDATA(121)",
	OutTemp       => APUFCMLOADDATA_OUT(121),
	Paths         => (0 => (CPMFCMCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => APUFCMLOADDATA(122),
	GlitchData    => APUFCMLOADDATA122_GlitchData,
	OutSignalName => "APUFCMLOADDATA(122)",
	OutTemp       => APUFCMLOADDATA_OUT(122),
	Paths         => (0 => (CPMFCMCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => APUFCMLOADDATA(123),
	GlitchData    => APUFCMLOADDATA123_GlitchData,
	OutSignalName => "APUFCMLOADDATA(123)",
	OutTemp       => APUFCMLOADDATA_OUT(123),
	Paths         => (0 => (CPMFCMCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => APUFCMLOADDATA(124),
	GlitchData    => APUFCMLOADDATA124_GlitchData,
	OutSignalName => "APUFCMLOADDATA(124)",
	OutTemp       => APUFCMLOADDATA_OUT(124),
	Paths         => (0 => (CPMFCMCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => APUFCMLOADDATA(125),
	GlitchData    => APUFCMLOADDATA125_GlitchData,
	OutSignalName => "APUFCMLOADDATA(125)",
	OutTemp       => APUFCMLOADDATA_OUT(125),
	Paths         => (0 => (CPMFCMCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => APUFCMLOADDATA(126),
	GlitchData    => APUFCMLOADDATA126_GlitchData,
	OutSignalName => "APUFCMLOADDATA(126)",
	OutTemp       => APUFCMLOADDATA_OUT(126),
	Paths         => (0 => (CPMFCMCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => APUFCMLOADDATA(127),
	GlitchData    => APUFCMLOADDATA127_GlitchData,
	OutSignalName => "APUFCMLOADDATA(127)",
	OutTemp       => APUFCMLOADDATA_OUT(127),
	Paths         => (0 => (CPMFCMCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => APUFCMLOADDVALID,
	GlitchData    => APUFCMLOADDVALID_GlitchData,
	OutSignalName => "APUFCMLOADDVALID",
	OutTemp       => APUFCMLOADDVALID_OUT,
	Paths         => (0 => (CPMFCMCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => APUFCMMSRFE0,
	GlitchData    => APUFCMMSRFE0_GlitchData,
	OutSignalName => "APUFCMMSRFE0",
	OutTemp       => APUFCMMSRFE0_OUT,
	Paths         => (0 => (CPMFCMCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => APUFCMMSRFE1,
	GlitchData    => APUFCMMSRFE1_GlitchData,
	OutSignalName => "APUFCMMSRFE1",
	OutTemp       => APUFCMMSRFE1_OUT,
	Paths         => (0 => (CPMFCMCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => APUFCMNEXTINSTRREADY,
	GlitchData    => APUFCMNEXTINSTRREADY_GlitchData,
	OutSignalName => "APUFCMNEXTINSTRREADY",
	OutTemp       => APUFCMNEXTINSTRREADY_OUT,
	Paths         => (0 => (CPMFCMCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => APUFCMOPERANDVALID,
	GlitchData    => APUFCMOPERANDVALID_GlitchData,
	OutSignalName => "APUFCMOPERANDVALID",
	OutTemp       => APUFCMOPERANDVALID_OUT,
	Paths         => (0 => (CPMFCMCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => APUFCMRADATA(0),
	GlitchData    => APUFCMRADATA0_GlitchData,
	OutSignalName => "APUFCMRADATA(0)",
	OutTemp       => APUFCMRADATA_OUT(0),
	Paths         => (0 => (CPMFCMCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => APUFCMRADATA(1),
	GlitchData    => APUFCMRADATA1_GlitchData,
	OutSignalName => "APUFCMRADATA(1)",
	OutTemp       => APUFCMRADATA_OUT(1),
	Paths         => (0 => (CPMFCMCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => APUFCMRADATA(2),
	GlitchData    => APUFCMRADATA2_GlitchData,
	OutSignalName => "APUFCMRADATA(2)",
	OutTemp       => APUFCMRADATA_OUT(2),
	Paths         => (0 => (CPMFCMCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => APUFCMRADATA(3),
	GlitchData    => APUFCMRADATA3_GlitchData,
	OutSignalName => "APUFCMRADATA(3)",
	OutTemp       => APUFCMRADATA_OUT(3),
	Paths         => (0 => (CPMFCMCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => APUFCMRADATA(4),
	GlitchData    => APUFCMRADATA4_GlitchData,
	OutSignalName => "APUFCMRADATA(4)",
	OutTemp       => APUFCMRADATA_OUT(4),
	Paths         => (0 => (CPMFCMCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => APUFCMRADATA(5),
	GlitchData    => APUFCMRADATA5_GlitchData,
	OutSignalName => "APUFCMRADATA(5)",
	OutTemp       => APUFCMRADATA_OUT(5),
	Paths         => (0 => (CPMFCMCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => APUFCMRADATA(6),
	GlitchData    => APUFCMRADATA6_GlitchData,
	OutSignalName => "APUFCMRADATA(6)",
	OutTemp       => APUFCMRADATA_OUT(6),
	Paths         => (0 => (CPMFCMCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => APUFCMRADATA(7),
	GlitchData    => APUFCMRADATA7_GlitchData,
	OutSignalName => "APUFCMRADATA(7)",
	OutTemp       => APUFCMRADATA_OUT(7),
	Paths         => (0 => (CPMFCMCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => APUFCMRADATA(8),
	GlitchData    => APUFCMRADATA8_GlitchData,
	OutSignalName => "APUFCMRADATA(8)",
	OutTemp       => APUFCMRADATA_OUT(8),
	Paths         => (0 => (CPMFCMCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => APUFCMRADATA(9),
	GlitchData    => APUFCMRADATA9_GlitchData,
	OutSignalName => "APUFCMRADATA(9)",
	OutTemp       => APUFCMRADATA_OUT(9),
	Paths         => (0 => (CPMFCMCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => APUFCMRADATA(10),
	GlitchData    => APUFCMRADATA10_GlitchData,
	OutSignalName => "APUFCMRADATA(10)",
	OutTemp       => APUFCMRADATA_OUT(10),
	Paths         => (0 => (CPMFCMCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => APUFCMRADATA(11),
	GlitchData    => APUFCMRADATA11_GlitchData,
	OutSignalName => "APUFCMRADATA(11)",
	OutTemp       => APUFCMRADATA_OUT(11),
	Paths         => (0 => (CPMFCMCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => APUFCMRADATA(12),
	GlitchData    => APUFCMRADATA12_GlitchData,
	OutSignalName => "APUFCMRADATA(12)",
	OutTemp       => APUFCMRADATA_OUT(12),
	Paths         => (0 => (CPMFCMCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => APUFCMRADATA(13),
	GlitchData    => APUFCMRADATA13_GlitchData,
	OutSignalName => "APUFCMRADATA(13)",
	OutTemp       => APUFCMRADATA_OUT(13),
	Paths         => (0 => (CPMFCMCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => APUFCMRADATA(14),
	GlitchData    => APUFCMRADATA14_GlitchData,
	OutSignalName => "APUFCMRADATA(14)",
	OutTemp       => APUFCMRADATA_OUT(14),
	Paths         => (0 => (CPMFCMCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => APUFCMRADATA(15),
	GlitchData    => APUFCMRADATA15_GlitchData,
	OutSignalName => "APUFCMRADATA(15)",
	OutTemp       => APUFCMRADATA_OUT(15),
	Paths         => (0 => (CPMFCMCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => APUFCMRADATA(16),
	GlitchData    => APUFCMRADATA16_GlitchData,
	OutSignalName => "APUFCMRADATA(16)",
	OutTemp       => APUFCMRADATA_OUT(16),
	Paths         => (0 => (CPMFCMCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => APUFCMRADATA(17),
	GlitchData    => APUFCMRADATA17_GlitchData,
	OutSignalName => "APUFCMRADATA(17)",
	OutTemp       => APUFCMRADATA_OUT(17),
	Paths         => (0 => (CPMFCMCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => APUFCMRADATA(18),
	GlitchData    => APUFCMRADATA18_GlitchData,
	OutSignalName => "APUFCMRADATA(18)",
	OutTemp       => APUFCMRADATA_OUT(18),
	Paths         => (0 => (CPMFCMCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => APUFCMRADATA(19),
	GlitchData    => APUFCMRADATA19_GlitchData,
	OutSignalName => "APUFCMRADATA(19)",
	OutTemp       => APUFCMRADATA_OUT(19),
	Paths         => (0 => (CPMFCMCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => APUFCMRADATA(20),
	GlitchData    => APUFCMRADATA20_GlitchData,
	OutSignalName => "APUFCMRADATA(20)",
	OutTemp       => APUFCMRADATA_OUT(20),
	Paths         => (0 => (CPMFCMCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => APUFCMRADATA(21),
	GlitchData    => APUFCMRADATA21_GlitchData,
	OutSignalName => "APUFCMRADATA(21)",
	OutTemp       => APUFCMRADATA_OUT(21),
	Paths         => (0 => (CPMFCMCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => APUFCMRADATA(22),
	GlitchData    => APUFCMRADATA22_GlitchData,
	OutSignalName => "APUFCMRADATA(22)",
	OutTemp       => APUFCMRADATA_OUT(22),
	Paths         => (0 => (CPMFCMCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => APUFCMRADATA(23),
	GlitchData    => APUFCMRADATA23_GlitchData,
	OutSignalName => "APUFCMRADATA(23)",
	OutTemp       => APUFCMRADATA_OUT(23),
	Paths         => (0 => (CPMFCMCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => APUFCMRADATA(24),
	GlitchData    => APUFCMRADATA24_GlitchData,
	OutSignalName => "APUFCMRADATA(24)",
	OutTemp       => APUFCMRADATA_OUT(24),
	Paths         => (0 => (CPMFCMCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => APUFCMRADATA(25),
	GlitchData    => APUFCMRADATA25_GlitchData,
	OutSignalName => "APUFCMRADATA(25)",
	OutTemp       => APUFCMRADATA_OUT(25),
	Paths         => (0 => (CPMFCMCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => APUFCMRADATA(26),
	GlitchData    => APUFCMRADATA26_GlitchData,
	OutSignalName => "APUFCMRADATA(26)",
	OutTemp       => APUFCMRADATA_OUT(26),
	Paths         => (0 => (CPMFCMCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => APUFCMRADATA(27),
	GlitchData    => APUFCMRADATA27_GlitchData,
	OutSignalName => "APUFCMRADATA(27)",
	OutTemp       => APUFCMRADATA_OUT(27),
	Paths         => (0 => (CPMFCMCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => APUFCMRADATA(28),
	GlitchData    => APUFCMRADATA28_GlitchData,
	OutSignalName => "APUFCMRADATA(28)",
	OutTemp       => APUFCMRADATA_OUT(28),
	Paths         => (0 => (CPMFCMCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => APUFCMRADATA(29),
	GlitchData    => APUFCMRADATA29_GlitchData,
	OutSignalName => "APUFCMRADATA(29)",
	OutTemp       => APUFCMRADATA_OUT(29),
	Paths         => (0 => (CPMFCMCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => APUFCMRADATA(30),
	GlitchData    => APUFCMRADATA30_GlitchData,
	OutSignalName => "APUFCMRADATA(30)",
	OutTemp       => APUFCMRADATA_OUT(30),
	Paths         => (0 => (CPMFCMCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => APUFCMRADATA(31),
	GlitchData    => APUFCMRADATA31_GlitchData,
	OutSignalName => "APUFCMRADATA(31)",
	OutTemp       => APUFCMRADATA_OUT(31),
	Paths         => (0 => (CPMFCMCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => APUFCMRBDATA(0),
	GlitchData    => APUFCMRBDATA0_GlitchData,
	OutSignalName => "APUFCMRBDATA(0)",
	OutTemp       => APUFCMRBDATA_OUT(0),
	Paths         => (0 => (CPMFCMCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => APUFCMRBDATA(1),
	GlitchData    => APUFCMRBDATA1_GlitchData,
	OutSignalName => "APUFCMRBDATA(1)",
	OutTemp       => APUFCMRBDATA_OUT(1),
	Paths         => (0 => (CPMFCMCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => APUFCMRBDATA(2),
	GlitchData    => APUFCMRBDATA2_GlitchData,
	OutSignalName => "APUFCMRBDATA(2)",
	OutTemp       => APUFCMRBDATA_OUT(2),
	Paths         => (0 => (CPMFCMCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => APUFCMRBDATA(3),
	GlitchData    => APUFCMRBDATA3_GlitchData,
	OutSignalName => "APUFCMRBDATA(3)",
	OutTemp       => APUFCMRBDATA_OUT(3),
	Paths         => (0 => (CPMFCMCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => APUFCMRBDATA(4),
	GlitchData    => APUFCMRBDATA4_GlitchData,
	OutSignalName => "APUFCMRBDATA(4)",
	OutTemp       => APUFCMRBDATA_OUT(4),
	Paths         => (0 => (CPMFCMCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => APUFCMRBDATA(5),
	GlitchData    => APUFCMRBDATA5_GlitchData,
	OutSignalName => "APUFCMRBDATA(5)",
	OutTemp       => APUFCMRBDATA_OUT(5),
	Paths         => (0 => (CPMFCMCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => APUFCMRBDATA(6),
	GlitchData    => APUFCMRBDATA6_GlitchData,
	OutSignalName => "APUFCMRBDATA(6)",
	OutTemp       => APUFCMRBDATA_OUT(6),
	Paths         => (0 => (CPMFCMCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => APUFCMRBDATA(7),
	GlitchData    => APUFCMRBDATA7_GlitchData,
	OutSignalName => "APUFCMRBDATA(7)",
	OutTemp       => APUFCMRBDATA_OUT(7),
	Paths         => (0 => (CPMFCMCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => APUFCMRBDATA(8),
	GlitchData    => APUFCMRBDATA8_GlitchData,
	OutSignalName => "APUFCMRBDATA(8)",
	OutTemp       => APUFCMRBDATA_OUT(8),
	Paths         => (0 => (CPMFCMCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => APUFCMRBDATA(9),
	GlitchData    => APUFCMRBDATA9_GlitchData,
	OutSignalName => "APUFCMRBDATA(9)",
	OutTemp       => APUFCMRBDATA_OUT(9),
	Paths         => (0 => (CPMFCMCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => APUFCMRBDATA(10),
	GlitchData    => APUFCMRBDATA10_GlitchData,
	OutSignalName => "APUFCMRBDATA(10)",
	OutTemp       => APUFCMRBDATA_OUT(10),
	Paths         => (0 => (CPMFCMCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => APUFCMRBDATA(11),
	GlitchData    => APUFCMRBDATA11_GlitchData,
	OutSignalName => "APUFCMRBDATA(11)",
	OutTemp       => APUFCMRBDATA_OUT(11),
	Paths         => (0 => (CPMFCMCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => APUFCMRBDATA(12),
	GlitchData    => APUFCMRBDATA12_GlitchData,
	OutSignalName => "APUFCMRBDATA(12)",
	OutTemp       => APUFCMRBDATA_OUT(12),
	Paths         => (0 => (CPMFCMCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => APUFCMRBDATA(13),
	GlitchData    => APUFCMRBDATA13_GlitchData,
	OutSignalName => "APUFCMRBDATA(13)",
	OutTemp       => APUFCMRBDATA_OUT(13),
	Paths         => (0 => (CPMFCMCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => APUFCMRBDATA(14),
	GlitchData    => APUFCMRBDATA14_GlitchData,
	OutSignalName => "APUFCMRBDATA(14)",
	OutTemp       => APUFCMRBDATA_OUT(14),
	Paths         => (0 => (CPMFCMCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => APUFCMRBDATA(15),
	GlitchData    => APUFCMRBDATA15_GlitchData,
	OutSignalName => "APUFCMRBDATA(15)",
	OutTemp       => APUFCMRBDATA_OUT(15),
	Paths         => (0 => (CPMFCMCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => APUFCMRBDATA(16),
	GlitchData    => APUFCMRBDATA16_GlitchData,
	OutSignalName => "APUFCMRBDATA(16)",
	OutTemp       => APUFCMRBDATA_OUT(16),
	Paths         => (0 => (CPMFCMCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => APUFCMRBDATA(17),
	GlitchData    => APUFCMRBDATA17_GlitchData,
	OutSignalName => "APUFCMRBDATA(17)",
	OutTemp       => APUFCMRBDATA_OUT(17),
	Paths         => (0 => (CPMFCMCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => APUFCMRBDATA(18),
	GlitchData    => APUFCMRBDATA18_GlitchData,
	OutSignalName => "APUFCMRBDATA(18)",
	OutTemp       => APUFCMRBDATA_OUT(18),
	Paths         => (0 => (CPMFCMCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => APUFCMRBDATA(19),
	GlitchData    => APUFCMRBDATA19_GlitchData,
	OutSignalName => "APUFCMRBDATA(19)",
	OutTemp       => APUFCMRBDATA_OUT(19),
	Paths         => (0 => (CPMFCMCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => APUFCMRBDATA(20),
	GlitchData    => APUFCMRBDATA20_GlitchData,
	OutSignalName => "APUFCMRBDATA(20)",
	OutTemp       => APUFCMRBDATA_OUT(20),
	Paths         => (0 => (CPMFCMCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => APUFCMRBDATA(21),
	GlitchData    => APUFCMRBDATA21_GlitchData,
	OutSignalName => "APUFCMRBDATA(21)",
	OutTemp       => APUFCMRBDATA_OUT(21),
	Paths         => (0 => (CPMFCMCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => APUFCMRBDATA(22),
	GlitchData    => APUFCMRBDATA22_GlitchData,
	OutSignalName => "APUFCMRBDATA(22)",
	OutTemp       => APUFCMRBDATA_OUT(22),
	Paths         => (0 => (CPMFCMCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => APUFCMRBDATA(23),
	GlitchData    => APUFCMRBDATA23_GlitchData,
	OutSignalName => "APUFCMRBDATA(23)",
	OutTemp       => APUFCMRBDATA_OUT(23),
	Paths         => (0 => (CPMFCMCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => APUFCMRBDATA(24),
	GlitchData    => APUFCMRBDATA24_GlitchData,
	OutSignalName => "APUFCMRBDATA(24)",
	OutTemp       => APUFCMRBDATA_OUT(24),
	Paths         => (0 => (CPMFCMCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => APUFCMRBDATA(25),
	GlitchData    => APUFCMRBDATA25_GlitchData,
	OutSignalName => "APUFCMRBDATA(25)",
	OutTemp       => APUFCMRBDATA_OUT(25),
	Paths         => (0 => (CPMFCMCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => APUFCMRBDATA(26),
	GlitchData    => APUFCMRBDATA26_GlitchData,
	OutSignalName => "APUFCMRBDATA(26)",
	OutTemp       => APUFCMRBDATA_OUT(26),
	Paths         => (0 => (CPMFCMCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => APUFCMRBDATA(27),
	GlitchData    => APUFCMRBDATA27_GlitchData,
	OutSignalName => "APUFCMRBDATA(27)",
	OutTemp       => APUFCMRBDATA_OUT(27),
	Paths         => (0 => (CPMFCMCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => APUFCMRBDATA(28),
	GlitchData    => APUFCMRBDATA28_GlitchData,
	OutSignalName => "APUFCMRBDATA(28)",
	OutTemp       => APUFCMRBDATA_OUT(28),
	Paths         => (0 => (CPMFCMCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => APUFCMRBDATA(29),
	GlitchData    => APUFCMRBDATA29_GlitchData,
	OutSignalName => "APUFCMRBDATA(29)",
	OutTemp       => APUFCMRBDATA_OUT(29),
	Paths         => (0 => (CPMFCMCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => APUFCMRBDATA(30),
	GlitchData    => APUFCMRBDATA30_GlitchData,
	OutSignalName => "APUFCMRBDATA(30)",
	OutTemp       => APUFCMRBDATA_OUT(30),
	Paths         => (0 => (CPMFCMCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => APUFCMRBDATA(31),
	GlitchData    => APUFCMRBDATA31_GlitchData,
	OutSignalName => "APUFCMRBDATA(31)",
	OutTemp       => APUFCMRBDATA_OUT(31),
	Paths         => (0 => (CPMFCMCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => APUFCMWRITEBACKOK,
	GlitchData    => APUFCMWRITEBACKOK_GlitchData,
	OutSignalName => "APUFCMWRITEBACKOK",
	OutTemp       => APUFCMWRITEBACKOK_OUT,
	Paths         => (0 => (CPMFCMCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => C440CPMCORESLEEPREQ,
	GlitchData    => C440CPMCORESLEEPREQ_GlitchData,
	OutSignalName => "C440CPMCORESLEEPREQ",
	OutTemp       => C440CPMCORESLEEPREQ_OUT,
	Paths         => (0 => (CPMC440CLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => C440CPMDECIRPTREQ,
	GlitchData    => C440CPMDECIRPTREQ_GlitchData,
	OutSignalName => "C440CPMDECIRPTREQ",
	OutTemp       => C440CPMDECIRPTREQ_OUT,
	Paths         => (0 => (CPMC440CLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => C440CPMFITIRPTREQ,
	GlitchData    => C440CPMFITIRPTREQ_GlitchData,
	OutSignalName => "C440CPMFITIRPTREQ",
	OutTemp       => C440CPMFITIRPTREQ_OUT,
	Paths         => (0 => (CPMC440CLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => C440CPMMSRCE,
	GlitchData    => C440CPMMSRCE_GlitchData,
	OutSignalName => "C440CPMMSRCE",
	OutTemp       => C440CPMMSRCE_OUT,
	Paths         => (0 => (CPMC440CLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => C440CPMMSREE,
	GlitchData    => C440CPMMSREE_GlitchData,
	OutSignalName => "C440CPMMSREE",
	OutTemp       => C440CPMMSREE_OUT,
	Paths         => (0 => (CPMC440CLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => C440CPMTIMERRESETREQ,
	GlitchData    => C440CPMTIMERRESETREQ_GlitchData,
	OutSignalName => "C440CPMTIMERRESETREQ",
	OutTemp       => C440CPMTIMERRESETREQ_OUT,
	Paths         => (0 => (CPMC440CLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => C440CPMWDIRPTREQ,
	GlitchData    => C440CPMWDIRPTREQ_GlitchData,
	OutSignalName => "C440CPMWDIRPTREQ",
	OutTemp       => C440CPMWDIRPTREQ_OUT,
	Paths         => (0 => (CPMC440CLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => C440DBGSYSTEMCONTROL(0),
	GlitchData    => C440DBGSYSTEMCONTROL0_GlitchData,
	OutSignalName => "C440DBGSYSTEMCONTROL(0)",
	OutTemp       => C440DBGSYSTEMCONTROL_OUT(0),
	Paths         => (0 => (CPMC440CLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => C440DBGSYSTEMCONTROL(1),
	GlitchData    => C440DBGSYSTEMCONTROL1_GlitchData,
	OutSignalName => "C440DBGSYSTEMCONTROL(1)",
	OutTemp       => C440DBGSYSTEMCONTROL_OUT(1),
	Paths         => (0 => (CPMC440CLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => C440DBGSYSTEMCONTROL(2),
	GlitchData    => C440DBGSYSTEMCONTROL2_GlitchData,
	OutSignalName => "C440DBGSYSTEMCONTROL(2)",
	OutTemp       => C440DBGSYSTEMCONTROL_OUT(2),
	Paths         => (0 => (CPMC440CLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => C440DBGSYSTEMCONTROL(3),
	GlitchData    => C440DBGSYSTEMCONTROL3_GlitchData,
	OutSignalName => "C440DBGSYSTEMCONTROL(3)",
	OutTemp       => C440DBGSYSTEMCONTROL_OUT(3),
	Paths         => (0 => (CPMC440CLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => C440DBGSYSTEMCONTROL(4),
	GlitchData    => C440DBGSYSTEMCONTROL4_GlitchData,
	OutSignalName => "C440DBGSYSTEMCONTROL(4)",
	OutTemp       => C440DBGSYSTEMCONTROL_OUT(4),
	Paths         => (0 => (CPMC440CLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => C440DBGSYSTEMCONTROL(5),
	GlitchData    => C440DBGSYSTEMCONTROL5_GlitchData,
	OutSignalName => "C440DBGSYSTEMCONTROL(5)",
	OutTemp       => C440DBGSYSTEMCONTROL_OUT(5),
	Paths         => (0 => (CPMC440CLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => C440DBGSYSTEMCONTROL(6),
	GlitchData    => C440DBGSYSTEMCONTROL6_GlitchData,
	OutSignalName => "C440DBGSYSTEMCONTROL(6)",
	OutTemp       => C440DBGSYSTEMCONTROL_OUT(6),
	Paths         => (0 => (CPMC440CLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => C440DBGSYSTEMCONTROL(7),
	GlitchData    => C440DBGSYSTEMCONTROL7_GlitchData,
	OutSignalName => "C440DBGSYSTEMCONTROL(7)",
	OutTemp       => C440DBGSYSTEMCONTROL_OUT(7),
	Paths         => (0 => (CPMC440CLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => C440JTGTDO,
	GlitchData    => C440JTGTDO_GlitchData,
	OutSignalName => "C440JTGTDO",
	OutTemp       => C440JTGTDO_OUT,
	Paths         => (0 => (JTGC440TCK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => C440JTGTDOEN,
	GlitchData    => C440JTGTDOEN_GlitchData,
	OutSignalName => "C440JTGTDOEN",
	OutTemp       => C440JTGTDOEN_OUT,
	Paths         => (0 => (JTGC440TCK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => C440MACHINECHECK,
	GlitchData    => C440MACHINECHECK_GlitchData,
	OutSignalName => "C440MACHINECHECK",
	OutTemp       => C440MACHINECHECK_OUT,
	Paths         => (0 => (CPMC440CLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => C440RSTCHIPRESETREQ,
	GlitchData    => C440RSTCHIPRESETREQ_GlitchData,
	OutSignalName => "C440RSTCHIPRESETREQ",
	OutTemp       => C440RSTCHIPRESETREQ_OUT,
	Paths         => (0 => (CPMINTERCONNECTCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => C440RSTCORERESETREQ,
	GlitchData    => C440RSTCORERESETREQ_GlitchData,
	OutSignalName => "C440RSTCORERESETREQ",
	OutTemp       => C440RSTCORERESETREQ_OUT,
	Paths         => (0 => (CPMINTERCONNECTCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => C440RSTSYSTEMRESETREQ,
	GlitchData    => C440RSTSYSTEMRESETREQ_GlitchData,
	OutSignalName => "C440RSTSYSTEMRESETREQ",
	OutTemp       => C440RSTSYSTEMRESETREQ_OUT,
	Paths         => (0 => (CPMINTERCONNECTCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => C440TRCBRANCHSTATUS(0),
	GlitchData    => C440TRCBRANCHSTATUS0_GlitchData,
	OutSignalName => "C440TRCBRANCHSTATUS(0)",
	OutTemp       => C440TRCBRANCHSTATUS_OUT(0),
	Paths         => (0 => (CPMC440CLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => C440TRCBRANCHSTATUS(1),
	GlitchData    => C440TRCBRANCHSTATUS1_GlitchData,
	OutSignalName => "C440TRCBRANCHSTATUS(1)",
	OutTemp       => C440TRCBRANCHSTATUS_OUT(1),
	Paths         => (0 => (CPMC440CLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => C440TRCBRANCHSTATUS(2),
	GlitchData    => C440TRCBRANCHSTATUS2_GlitchData,
	OutSignalName => "C440TRCBRANCHSTATUS(2)",
	OutTemp       => C440TRCBRANCHSTATUS_OUT(2),
	Paths         => (0 => (CPMC440CLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => C440TRCCYCLE,
	GlitchData    => C440TRCCYCLE_GlitchData,
	OutSignalName => "C440TRCCYCLE",
	OutTemp       => C440TRCCYCLE_OUT,
	Paths         => (0 => (CPMC440CLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => C440TRCEXECUTIONSTATUS(0),
	GlitchData    => C440TRCEXECUTIONSTATUS0_GlitchData,
	OutSignalName => "C440TRCEXECUTIONSTATUS(0)",
	OutTemp       => C440TRCEXECUTIONSTATUS_OUT(0),
	Paths         => (0 => (CPMC440CLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => C440TRCEXECUTIONSTATUS(1),
	GlitchData    => C440TRCEXECUTIONSTATUS1_GlitchData,
	OutSignalName => "C440TRCEXECUTIONSTATUS(1)",
	OutTemp       => C440TRCEXECUTIONSTATUS_OUT(1),
	Paths         => (0 => (CPMC440CLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => C440TRCEXECUTIONSTATUS(2),
	GlitchData    => C440TRCEXECUTIONSTATUS2_GlitchData,
	OutSignalName => "C440TRCEXECUTIONSTATUS(2)",
	OutTemp       => C440TRCEXECUTIONSTATUS_OUT(2),
	Paths         => (0 => (CPMC440CLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => C440TRCEXECUTIONSTATUS(3),
	GlitchData    => C440TRCEXECUTIONSTATUS3_GlitchData,
	OutSignalName => "C440TRCEXECUTIONSTATUS(3)",
	OutTemp       => C440TRCEXECUTIONSTATUS_OUT(3),
	Paths         => (0 => (CPMC440CLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => C440TRCEXECUTIONSTATUS(4),
	GlitchData    => C440TRCEXECUTIONSTATUS4_GlitchData,
	OutSignalName => "C440TRCEXECUTIONSTATUS(4)",
	OutTemp       => C440TRCEXECUTIONSTATUS_OUT(4),
	Paths         => (0 => (CPMC440CLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => C440TRCTRACESTATUS(0),
	GlitchData    => C440TRCTRACESTATUS0_GlitchData,
	OutSignalName => "C440TRCTRACESTATUS(0)",
	OutTemp       => C440TRCTRACESTATUS_OUT(0),
	Paths         => (0 => (CPMC440CLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => C440TRCTRACESTATUS(1),
	GlitchData    => C440TRCTRACESTATUS1_GlitchData,
	OutSignalName => "C440TRCTRACESTATUS(1)",
	OutTemp       => C440TRCTRACESTATUS_OUT(1),
	Paths         => (0 => (CPMC440CLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => C440TRCTRACESTATUS(2),
	GlitchData    => C440TRCTRACESTATUS2_GlitchData,
	OutSignalName => "C440TRCTRACESTATUS(2)",
	OutTemp       => C440TRCTRACESTATUS_OUT(2),
	Paths         => (0 => (CPMC440CLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => C440TRCTRACESTATUS(3),
	GlitchData    => C440TRCTRACESTATUS3_GlitchData,
	OutSignalName => "C440TRCTRACESTATUS(3)",
	OutTemp       => C440TRCTRACESTATUS_OUT(3),
	Paths         => (0 => (CPMC440CLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => C440TRCTRACESTATUS(4),
	GlitchData    => C440TRCTRACESTATUS4_GlitchData,
	OutSignalName => "C440TRCTRACESTATUS(4)",
	OutTemp       => C440TRCTRACESTATUS_OUT(4),
	Paths         => (0 => (CPMC440CLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => C440TRCTRACESTATUS(5),
	GlitchData    => C440TRCTRACESTATUS5_GlitchData,
	OutSignalName => "C440TRCTRACESTATUS(5)",
	OutTemp       => C440TRCTRACESTATUS_OUT(5),
	Paths         => (0 => (CPMC440CLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => C440TRCTRACESTATUS(6),
	GlitchData    => C440TRCTRACESTATUS6_GlitchData,
	OutSignalName => "C440TRCTRACESTATUS(6)",
	OutTemp       => C440TRCTRACESTATUS_OUT(6),
	Paths         => (0 => (CPMC440CLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => C440TRCTRIGGEREVENTOUT,
	GlitchData    => C440TRCTRIGGEREVENTOUT_GlitchData,
	OutSignalName => "C440TRCTRIGGEREVENTOUT",
	OutTemp       => C440TRCTRIGGEREVENTOUT_OUT,
	Paths         => (0 => (CPMC440CLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => C440TRCTRIGGEREVENTTYPE(0),
	GlitchData    => C440TRCTRIGGEREVENTTYPE0_GlitchData,
	OutSignalName => "C440TRCTRIGGEREVENTTYPE(0)",
	OutTemp       => C440TRCTRIGGEREVENTTYPE_OUT(0),
	Paths         => (0 => (CPMC440CLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => C440TRCTRIGGEREVENTTYPE(1),
	GlitchData    => C440TRCTRIGGEREVENTTYPE1_GlitchData,
	OutSignalName => "C440TRCTRIGGEREVENTTYPE(1)",
	OutTemp       => C440TRCTRIGGEREVENTTYPE_OUT(1),
	Paths         => (0 => (CPMC440CLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => C440TRCTRIGGEREVENTTYPE(2),
	GlitchData    => C440TRCTRIGGEREVENTTYPE2_GlitchData,
	OutSignalName => "C440TRCTRIGGEREVENTTYPE(2)",
	OutTemp       => C440TRCTRIGGEREVENTTYPE_OUT(2),
	Paths         => (0 => (CPMC440CLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => C440TRCTRIGGEREVENTTYPE(3),
	GlitchData    => C440TRCTRIGGEREVENTTYPE3_GlitchData,
	OutSignalName => "C440TRCTRIGGEREVENTTYPE(3)",
	OutTemp       => C440TRCTRIGGEREVENTTYPE_OUT(3),
	Paths         => (0 => (CPMC440CLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => C440TRCTRIGGEREVENTTYPE(4),
	GlitchData    => C440TRCTRIGGEREVENTTYPE4_GlitchData,
	OutSignalName => "C440TRCTRIGGEREVENTTYPE(4)",
	OutTemp       => C440TRCTRIGGEREVENTTYPE_OUT(4),
	Paths         => (0 => (CPMC440CLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => C440TRCTRIGGEREVENTTYPE(5),
	GlitchData    => C440TRCTRIGGEREVENTTYPE5_GlitchData,
	OutSignalName => "C440TRCTRIGGEREVENTTYPE(5)",
	OutTemp       => C440TRCTRIGGEREVENTTYPE_OUT(5),
	Paths         => (0 => (CPMC440CLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => C440TRCTRIGGEREVENTTYPE(6),
	GlitchData    => C440TRCTRIGGEREVENTTYPE6_GlitchData,
	OutSignalName => "C440TRCTRIGGEREVENTTYPE(6)",
	OutTemp       => C440TRCTRIGGEREVENTTYPE_OUT(6),
	Paths         => (0 => (CPMC440CLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => C440TRCTRIGGEREVENTTYPE(7),
	GlitchData    => C440TRCTRIGGEREVENTTYPE7_GlitchData,
	OutSignalName => "C440TRCTRIGGEREVENTTYPE(7)",
	OutTemp       => C440TRCTRIGGEREVENTTYPE_OUT(7),
	Paths         => (0 => (CPMC440CLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => C440TRCTRIGGEREVENTTYPE(8),
	GlitchData    => C440TRCTRIGGEREVENTTYPE8_GlitchData,
	OutSignalName => "C440TRCTRIGGEREVENTTYPE(8)",
	OutTemp       => C440TRCTRIGGEREVENTTYPE_OUT(8),
	Paths         => (0 => (CPMC440CLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => C440TRCTRIGGEREVENTTYPE(9),
	GlitchData    => C440TRCTRIGGEREVENTTYPE9_GlitchData,
	OutSignalName => "C440TRCTRIGGEREVENTTYPE(9)",
	OutTemp       => C440TRCTRIGGEREVENTTYPE_OUT(9),
	Paths         => (0 => (CPMC440CLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => C440TRCTRIGGEREVENTTYPE(10),
	GlitchData    => C440TRCTRIGGEREVENTTYPE10_GlitchData,
	OutSignalName => "C440TRCTRIGGEREVENTTYPE(10)",
	OutTemp       => C440TRCTRIGGEREVENTTYPE_OUT(10),
	Paths         => (0 => (CPMC440CLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => C440TRCTRIGGEREVENTTYPE(11),
	GlitchData    => C440TRCTRIGGEREVENTTYPE11_GlitchData,
	OutSignalName => "C440TRCTRIGGEREVENTTYPE(11)",
	OutTemp       => C440TRCTRIGGEREVENTTYPE_OUT(11),
	Paths         => (0 => (CPMC440CLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => C440TRCTRIGGEREVENTTYPE(12),
	GlitchData    => C440TRCTRIGGEREVENTTYPE12_GlitchData,
	OutSignalName => "C440TRCTRIGGEREVENTTYPE(12)",
	OutTemp       => C440TRCTRIGGEREVENTTYPE_OUT(12),
	Paths         => (0 => (CPMC440CLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => C440TRCTRIGGEREVENTTYPE(13),
	GlitchData    => C440TRCTRIGGEREVENTTYPE13_GlitchData,
	OutSignalName => "C440TRCTRIGGEREVENTTYPE(13)",
	OutTemp       => C440TRCTRIGGEREVENTTYPE_OUT(13),
	Paths         => (0 => (CPMC440CLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => MIMCADDRESS(0),
	GlitchData    => MIMCADDRESS0_GlitchData,
	OutSignalName => "MIMCADDRESS(0)",
	OutTemp       => MIMCADDRESS_OUT(0),
	Paths         => (0 => (CPMMCCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => MIMCADDRESS(1),
	GlitchData    => MIMCADDRESS1_GlitchData,
	OutSignalName => "MIMCADDRESS(1)",
	OutTemp       => MIMCADDRESS_OUT(1),
	Paths         => (0 => (CPMMCCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => MIMCADDRESS(2),
	GlitchData    => MIMCADDRESS2_GlitchData,
	OutSignalName => "MIMCADDRESS(2)",
	OutTemp       => MIMCADDRESS_OUT(2),
	Paths         => (0 => (CPMMCCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => MIMCADDRESS(3),
	GlitchData    => MIMCADDRESS3_GlitchData,
	OutSignalName => "MIMCADDRESS(3)",
	OutTemp       => MIMCADDRESS_OUT(3),
	Paths         => (0 => (CPMMCCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => MIMCADDRESS(4),
	GlitchData    => MIMCADDRESS4_GlitchData,
	OutSignalName => "MIMCADDRESS(4)",
	OutTemp       => MIMCADDRESS_OUT(4),
	Paths         => (0 => (CPMMCCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => MIMCADDRESS(5),
	GlitchData    => MIMCADDRESS5_GlitchData,
	OutSignalName => "MIMCADDRESS(5)",
	OutTemp       => MIMCADDRESS_OUT(5),
	Paths         => (0 => (CPMMCCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => MIMCADDRESS(6),
	GlitchData    => MIMCADDRESS6_GlitchData,
	OutSignalName => "MIMCADDRESS(6)",
	OutTemp       => MIMCADDRESS_OUT(6),
	Paths         => (0 => (CPMMCCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => MIMCADDRESS(7),
	GlitchData    => MIMCADDRESS7_GlitchData,
	OutSignalName => "MIMCADDRESS(7)",
	OutTemp       => MIMCADDRESS_OUT(7),
	Paths         => (0 => (CPMMCCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => MIMCADDRESS(8),
	GlitchData    => MIMCADDRESS8_GlitchData,
	OutSignalName => "MIMCADDRESS(8)",
	OutTemp       => MIMCADDRESS_OUT(8),
	Paths         => (0 => (CPMMCCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => MIMCADDRESS(9),
	GlitchData    => MIMCADDRESS9_GlitchData,
	OutSignalName => "MIMCADDRESS(9)",
	OutTemp       => MIMCADDRESS_OUT(9),
	Paths         => (0 => (CPMMCCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => MIMCADDRESS(10),
	GlitchData    => MIMCADDRESS10_GlitchData,
	OutSignalName => "MIMCADDRESS(10)",
	OutTemp       => MIMCADDRESS_OUT(10),
	Paths         => (0 => (CPMMCCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => MIMCADDRESS(11),
	GlitchData    => MIMCADDRESS11_GlitchData,
	OutSignalName => "MIMCADDRESS(11)",
	OutTemp       => MIMCADDRESS_OUT(11),
	Paths         => (0 => (CPMMCCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => MIMCADDRESS(12),
	GlitchData    => MIMCADDRESS12_GlitchData,
	OutSignalName => "MIMCADDRESS(12)",
	OutTemp       => MIMCADDRESS_OUT(12),
	Paths         => (0 => (CPMMCCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => MIMCADDRESS(13),
	GlitchData    => MIMCADDRESS13_GlitchData,
	OutSignalName => "MIMCADDRESS(13)",
	OutTemp       => MIMCADDRESS_OUT(13),
	Paths         => (0 => (CPMMCCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => MIMCADDRESS(14),
	GlitchData    => MIMCADDRESS14_GlitchData,
	OutSignalName => "MIMCADDRESS(14)",
	OutTemp       => MIMCADDRESS_OUT(14),
	Paths         => (0 => (CPMMCCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => MIMCADDRESS(15),
	GlitchData    => MIMCADDRESS15_GlitchData,
	OutSignalName => "MIMCADDRESS(15)",
	OutTemp       => MIMCADDRESS_OUT(15),
	Paths         => (0 => (CPMMCCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => MIMCADDRESS(16),
	GlitchData    => MIMCADDRESS16_GlitchData,
	OutSignalName => "MIMCADDRESS(16)",
	OutTemp       => MIMCADDRESS_OUT(16),
	Paths         => (0 => (CPMMCCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => MIMCADDRESS(17),
	GlitchData    => MIMCADDRESS17_GlitchData,
	OutSignalName => "MIMCADDRESS(17)",
	OutTemp       => MIMCADDRESS_OUT(17),
	Paths         => (0 => (CPMMCCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => MIMCADDRESS(18),
	GlitchData    => MIMCADDRESS18_GlitchData,
	OutSignalName => "MIMCADDRESS(18)",
	OutTemp       => MIMCADDRESS_OUT(18),
	Paths         => (0 => (CPMMCCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => MIMCADDRESS(19),
	GlitchData    => MIMCADDRESS19_GlitchData,
	OutSignalName => "MIMCADDRESS(19)",
	OutTemp       => MIMCADDRESS_OUT(19),
	Paths         => (0 => (CPMMCCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => MIMCADDRESS(20),
	GlitchData    => MIMCADDRESS20_GlitchData,
	OutSignalName => "MIMCADDRESS(20)",
	OutTemp       => MIMCADDRESS_OUT(20),
	Paths         => (0 => (CPMMCCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => MIMCADDRESS(21),
	GlitchData    => MIMCADDRESS21_GlitchData,
	OutSignalName => "MIMCADDRESS(21)",
	OutTemp       => MIMCADDRESS_OUT(21),
	Paths         => (0 => (CPMMCCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => MIMCADDRESS(22),
	GlitchData    => MIMCADDRESS22_GlitchData,
	OutSignalName => "MIMCADDRESS(22)",
	OutTemp       => MIMCADDRESS_OUT(22),
	Paths         => (0 => (CPMMCCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => MIMCADDRESS(23),
	GlitchData    => MIMCADDRESS23_GlitchData,
	OutSignalName => "MIMCADDRESS(23)",
	OutTemp       => MIMCADDRESS_OUT(23),
	Paths         => (0 => (CPMMCCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => MIMCADDRESS(24),
	GlitchData    => MIMCADDRESS24_GlitchData,
	OutSignalName => "MIMCADDRESS(24)",
	OutTemp       => MIMCADDRESS_OUT(24),
	Paths         => (0 => (CPMMCCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => MIMCADDRESS(25),
	GlitchData    => MIMCADDRESS25_GlitchData,
	OutSignalName => "MIMCADDRESS(25)",
	OutTemp       => MIMCADDRESS_OUT(25),
	Paths         => (0 => (CPMMCCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => MIMCADDRESS(26),
	GlitchData    => MIMCADDRESS26_GlitchData,
	OutSignalName => "MIMCADDRESS(26)",
	OutTemp       => MIMCADDRESS_OUT(26),
	Paths         => (0 => (CPMMCCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => MIMCADDRESS(27),
	GlitchData    => MIMCADDRESS27_GlitchData,
	OutSignalName => "MIMCADDRESS(27)",
	OutTemp       => MIMCADDRESS_OUT(27),
	Paths         => (0 => (CPMMCCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => MIMCADDRESS(28),
	GlitchData    => MIMCADDRESS28_GlitchData,
	OutSignalName => "MIMCADDRESS(28)",
	OutTemp       => MIMCADDRESS_OUT(28),
	Paths         => (0 => (CPMMCCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => MIMCADDRESS(29),
	GlitchData    => MIMCADDRESS29_GlitchData,
	OutSignalName => "MIMCADDRESS(29)",
	OutTemp       => MIMCADDRESS_OUT(29),
	Paths         => (0 => (CPMMCCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => MIMCADDRESS(30),
	GlitchData    => MIMCADDRESS30_GlitchData,
	OutSignalName => "MIMCADDRESS(30)",
	OutTemp       => MIMCADDRESS_OUT(30),
	Paths         => (0 => (CPMMCCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => MIMCADDRESS(31),
	GlitchData    => MIMCADDRESS31_GlitchData,
	OutSignalName => "MIMCADDRESS(31)",
	OutTemp       => MIMCADDRESS_OUT(31),
	Paths         => (0 => (CPMMCCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => MIMCADDRESS(32),
	GlitchData    => MIMCADDRESS32_GlitchData,
	OutSignalName => "MIMCADDRESS(32)",
	OutTemp       => MIMCADDRESS_OUT(32),
	Paths         => (0 => (CPMMCCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => MIMCADDRESS(33),
	GlitchData    => MIMCADDRESS33_GlitchData,
	OutSignalName => "MIMCADDRESS(33)",
	OutTemp       => MIMCADDRESS_OUT(33),
	Paths         => (0 => (CPMMCCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => MIMCADDRESS(34),
	GlitchData    => MIMCADDRESS34_GlitchData,
	OutSignalName => "MIMCADDRESS(34)",
	OutTemp       => MIMCADDRESS_OUT(34),
	Paths         => (0 => (CPMMCCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => MIMCADDRESS(35),
	GlitchData    => MIMCADDRESS35_GlitchData,
	OutSignalName => "MIMCADDRESS(35)",
	OutTemp       => MIMCADDRESS_OUT(35),
	Paths         => (0 => (CPMMCCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => MIMCADDRESSVALID,
	GlitchData    => MIMCADDRESSVALID_GlitchData,
	OutSignalName => "MIMCADDRESSVALID",
	OutTemp       => MIMCADDRESSVALID_OUT,
	Paths         => (0 => (CPMMCCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => MIMCBANKCONFLICT,
	GlitchData    => MIMCBANKCONFLICT_GlitchData,
	OutSignalName => "MIMCBANKCONFLICT",
	OutTemp       => MIMCBANKCONFLICT_OUT,
	Paths         => (0 => (CPMMCCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => MIMCBYTEENABLE(0),
	GlitchData    => MIMCBYTEENABLE0_GlitchData,
	OutSignalName => "MIMCBYTEENABLE(0)",
	OutTemp       => MIMCBYTEENABLE_OUT(0),
	Paths         => (0 => (CPMMCCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => MIMCBYTEENABLE(1),
	GlitchData    => MIMCBYTEENABLE1_GlitchData,
	OutSignalName => "MIMCBYTEENABLE(1)",
	OutTemp       => MIMCBYTEENABLE_OUT(1),
	Paths         => (0 => (CPMMCCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => MIMCBYTEENABLE(2),
	GlitchData    => MIMCBYTEENABLE2_GlitchData,
	OutSignalName => "MIMCBYTEENABLE(2)",
	OutTemp       => MIMCBYTEENABLE_OUT(2),
	Paths         => (0 => (CPMMCCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => MIMCBYTEENABLE(3),
	GlitchData    => MIMCBYTEENABLE3_GlitchData,
	OutSignalName => "MIMCBYTEENABLE(3)",
	OutTemp       => MIMCBYTEENABLE_OUT(3),
	Paths         => (0 => (CPMMCCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => MIMCBYTEENABLE(4),
	GlitchData    => MIMCBYTEENABLE4_GlitchData,
	OutSignalName => "MIMCBYTEENABLE(4)",
	OutTemp       => MIMCBYTEENABLE_OUT(4),
	Paths         => (0 => (CPMMCCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => MIMCBYTEENABLE(5),
	GlitchData    => MIMCBYTEENABLE5_GlitchData,
	OutSignalName => "MIMCBYTEENABLE(5)",
	OutTemp       => MIMCBYTEENABLE_OUT(5),
	Paths         => (0 => (CPMMCCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => MIMCBYTEENABLE(6),
	GlitchData    => MIMCBYTEENABLE6_GlitchData,
	OutSignalName => "MIMCBYTEENABLE(6)",
	OutTemp       => MIMCBYTEENABLE_OUT(6),
	Paths         => (0 => (CPMMCCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => MIMCBYTEENABLE(7),
	GlitchData    => MIMCBYTEENABLE7_GlitchData,
	OutSignalName => "MIMCBYTEENABLE(7)",
	OutTemp       => MIMCBYTEENABLE_OUT(7),
	Paths         => (0 => (CPMMCCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => MIMCBYTEENABLE(8),
	GlitchData    => MIMCBYTEENABLE8_GlitchData,
	OutSignalName => "MIMCBYTEENABLE(8)",
	OutTemp       => MIMCBYTEENABLE_OUT(8),
	Paths         => (0 => (CPMMCCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => MIMCBYTEENABLE(9),
	GlitchData    => MIMCBYTEENABLE9_GlitchData,
	OutSignalName => "MIMCBYTEENABLE(9)",
	OutTemp       => MIMCBYTEENABLE_OUT(9),
	Paths         => (0 => (CPMMCCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => MIMCBYTEENABLE(10),
	GlitchData    => MIMCBYTEENABLE10_GlitchData,
	OutSignalName => "MIMCBYTEENABLE(10)",
	OutTemp       => MIMCBYTEENABLE_OUT(10),
	Paths         => (0 => (CPMMCCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => MIMCBYTEENABLE(11),
	GlitchData    => MIMCBYTEENABLE11_GlitchData,
	OutSignalName => "MIMCBYTEENABLE(11)",
	OutTemp       => MIMCBYTEENABLE_OUT(11),
	Paths         => (0 => (CPMMCCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => MIMCBYTEENABLE(12),
	GlitchData    => MIMCBYTEENABLE12_GlitchData,
	OutSignalName => "MIMCBYTEENABLE(12)",
	OutTemp       => MIMCBYTEENABLE_OUT(12),
	Paths         => (0 => (CPMMCCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => MIMCBYTEENABLE(13),
	GlitchData    => MIMCBYTEENABLE13_GlitchData,
	OutSignalName => "MIMCBYTEENABLE(13)",
	OutTemp       => MIMCBYTEENABLE_OUT(13),
	Paths         => (0 => (CPMMCCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => MIMCBYTEENABLE(14),
	GlitchData    => MIMCBYTEENABLE14_GlitchData,
	OutSignalName => "MIMCBYTEENABLE(14)",
	OutTemp       => MIMCBYTEENABLE_OUT(14),
	Paths         => (0 => (CPMMCCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => MIMCBYTEENABLE(15),
	GlitchData    => MIMCBYTEENABLE15_GlitchData,
	OutSignalName => "MIMCBYTEENABLE(15)",
	OutTemp       => MIMCBYTEENABLE_OUT(15),
	Paths         => (0 => (CPMMCCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => MIMCREADNOTWRITE,
	GlitchData    => MIMCREADNOTWRITE_GlitchData,
	OutSignalName => "MIMCREADNOTWRITE",
	OutTemp       => MIMCREADNOTWRITE_OUT,
	Paths         => (0 => (CPMMCCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => MIMCROWCONFLICT,
	GlitchData    => MIMCROWCONFLICT_GlitchData,
	OutSignalName => "MIMCROWCONFLICT",
	OutTemp       => MIMCROWCONFLICT_OUT,
	Paths         => (0 => (CPMMCCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => MIMCWRITEDATA(0),
	GlitchData    => MIMCWRITEDATA0_GlitchData,
	OutSignalName => "MIMCWRITEDATA(0)",
	OutTemp       => MIMCWRITEDATA_OUT(0),
	Paths         => (0 => (CPMMCCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => MIMCWRITEDATA(1),
	GlitchData    => MIMCWRITEDATA1_GlitchData,
	OutSignalName => "MIMCWRITEDATA(1)",
	OutTemp       => MIMCWRITEDATA_OUT(1),
	Paths         => (0 => (CPMMCCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => MIMCWRITEDATA(2),
	GlitchData    => MIMCWRITEDATA2_GlitchData,
	OutSignalName => "MIMCWRITEDATA(2)",
	OutTemp       => MIMCWRITEDATA_OUT(2),
	Paths         => (0 => (CPMMCCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => MIMCWRITEDATA(3),
	GlitchData    => MIMCWRITEDATA3_GlitchData,
	OutSignalName => "MIMCWRITEDATA(3)",
	OutTemp       => MIMCWRITEDATA_OUT(3),
	Paths         => (0 => (CPMMCCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => MIMCWRITEDATA(4),
	GlitchData    => MIMCWRITEDATA4_GlitchData,
	OutSignalName => "MIMCWRITEDATA(4)",
	OutTemp       => MIMCWRITEDATA_OUT(4),
	Paths         => (0 => (CPMMCCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => MIMCWRITEDATA(5),
	GlitchData    => MIMCWRITEDATA5_GlitchData,
	OutSignalName => "MIMCWRITEDATA(5)",
	OutTemp       => MIMCWRITEDATA_OUT(5),
	Paths         => (0 => (CPMMCCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => MIMCWRITEDATA(6),
	GlitchData    => MIMCWRITEDATA6_GlitchData,
	OutSignalName => "MIMCWRITEDATA(6)",
	OutTemp       => MIMCWRITEDATA_OUT(6),
	Paths         => (0 => (CPMMCCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => MIMCWRITEDATA(7),
	GlitchData    => MIMCWRITEDATA7_GlitchData,
	OutSignalName => "MIMCWRITEDATA(7)",
	OutTemp       => MIMCWRITEDATA_OUT(7),
	Paths         => (0 => (CPMMCCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => MIMCWRITEDATA(8),
	GlitchData    => MIMCWRITEDATA8_GlitchData,
	OutSignalName => "MIMCWRITEDATA(8)",
	OutTemp       => MIMCWRITEDATA_OUT(8),
	Paths         => (0 => (CPMMCCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => MIMCWRITEDATA(9),
	GlitchData    => MIMCWRITEDATA9_GlitchData,
	OutSignalName => "MIMCWRITEDATA(9)",
	OutTemp       => MIMCWRITEDATA_OUT(9),
	Paths         => (0 => (CPMMCCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => MIMCWRITEDATA(10),
	GlitchData    => MIMCWRITEDATA10_GlitchData,
	OutSignalName => "MIMCWRITEDATA(10)",
	OutTemp       => MIMCWRITEDATA_OUT(10),
	Paths         => (0 => (CPMMCCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => MIMCWRITEDATA(11),
	GlitchData    => MIMCWRITEDATA11_GlitchData,
	OutSignalName => "MIMCWRITEDATA(11)",
	OutTemp       => MIMCWRITEDATA_OUT(11),
	Paths         => (0 => (CPMMCCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => MIMCWRITEDATA(12),
	GlitchData    => MIMCWRITEDATA12_GlitchData,
	OutSignalName => "MIMCWRITEDATA(12)",
	OutTemp       => MIMCWRITEDATA_OUT(12),
	Paths         => (0 => (CPMMCCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => MIMCWRITEDATA(13),
	GlitchData    => MIMCWRITEDATA13_GlitchData,
	OutSignalName => "MIMCWRITEDATA(13)",
	OutTemp       => MIMCWRITEDATA_OUT(13),
	Paths         => (0 => (CPMMCCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => MIMCWRITEDATA(14),
	GlitchData    => MIMCWRITEDATA14_GlitchData,
	OutSignalName => "MIMCWRITEDATA(14)",
	OutTemp       => MIMCWRITEDATA_OUT(14),
	Paths         => (0 => (CPMMCCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => MIMCWRITEDATA(15),
	GlitchData    => MIMCWRITEDATA15_GlitchData,
	OutSignalName => "MIMCWRITEDATA(15)",
	OutTemp       => MIMCWRITEDATA_OUT(15),
	Paths         => (0 => (CPMMCCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => MIMCWRITEDATA(16),
	GlitchData    => MIMCWRITEDATA16_GlitchData,
	OutSignalName => "MIMCWRITEDATA(16)",
	OutTemp       => MIMCWRITEDATA_OUT(16),
	Paths         => (0 => (CPMMCCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => MIMCWRITEDATA(17),
	GlitchData    => MIMCWRITEDATA17_GlitchData,
	OutSignalName => "MIMCWRITEDATA(17)",
	OutTemp       => MIMCWRITEDATA_OUT(17),
	Paths         => (0 => (CPMMCCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => MIMCWRITEDATA(18),
	GlitchData    => MIMCWRITEDATA18_GlitchData,
	OutSignalName => "MIMCWRITEDATA(18)",
	OutTemp       => MIMCWRITEDATA_OUT(18),
	Paths         => (0 => (CPMMCCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => MIMCWRITEDATA(19),
	GlitchData    => MIMCWRITEDATA19_GlitchData,
	OutSignalName => "MIMCWRITEDATA(19)",
	OutTemp       => MIMCWRITEDATA_OUT(19),
	Paths         => (0 => (CPMMCCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => MIMCWRITEDATA(20),
	GlitchData    => MIMCWRITEDATA20_GlitchData,
	OutSignalName => "MIMCWRITEDATA(20)",
	OutTemp       => MIMCWRITEDATA_OUT(20),
	Paths         => (0 => (CPMMCCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => MIMCWRITEDATA(21),
	GlitchData    => MIMCWRITEDATA21_GlitchData,
	OutSignalName => "MIMCWRITEDATA(21)",
	OutTemp       => MIMCWRITEDATA_OUT(21),
	Paths         => (0 => (CPMMCCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => MIMCWRITEDATA(22),
	GlitchData    => MIMCWRITEDATA22_GlitchData,
	OutSignalName => "MIMCWRITEDATA(22)",
	OutTemp       => MIMCWRITEDATA_OUT(22),
	Paths         => (0 => (CPMMCCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => MIMCWRITEDATA(23),
	GlitchData    => MIMCWRITEDATA23_GlitchData,
	OutSignalName => "MIMCWRITEDATA(23)",
	OutTemp       => MIMCWRITEDATA_OUT(23),
	Paths         => (0 => (CPMMCCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => MIMCWRITEDATA(24),
	GlitchData    => MIMCWRITEDATA24_GlitchData,
	OutSignalName => "MIMCWRITEDATA(24)",
	OutTemp       => MIMCWRITEDATA_OUT(24),
	Paths         => (0 => (CPMMCCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => MIMCWRITEDATA(25),
	GlitchData    => MIMCWRITEDATA25_GlitchData,
	OutSignalName => "MIMCWRITEDATA(25)",
	OutTemp       => MIMCWRITEDATA_OUT(25),
	Paths         => (0 => (CPMMCCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => MIMCWRITEDATA(26),
	GlitchData    => MIMCWRITEDATA26_GlitchData,
	OutSignalName => "MIMCWRITEDATA(26)",
	OutTemp       => MIMCWRITEDATA_OUT(26),
	Paths         => (0 => (CPMMCCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => MIMCWRITEDATA(27),
	GlitchData    => MIMCWRITEDATA27_GlitchData,
	OutSignalName => "MIMCWRITEDATA(27)",
	OutTemp       => MIMCWRITEDATA_OUT(27),
	Paths         => (0 => (CPMMCCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => MIMCWRITEDATA(28),
	GlitchData    => MIMCWRITEDATA28_GlitchData,
	OutSignalName => "MIMCWRITEDATA(28)",
	OutTemp       => MIMCWRITEDATA_OUT(28),
	Paths         => (0 => (CPMMCCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => MIMCWRITEDATA(29),
	GlitchData    => MIMCWRITEDATA29_GlitchData,
	OutSignalName => "MIMCWRITEDATA(29)",
	OutTemp       => MIMCWRITEDATA_OUT(29),
	Paths         => (0 => (CPMMCCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => MIMCWRITEDATA(30),
	GlitchData    => MIMCWRITEDATA30_GlitchData,
	OutSignalName => "MIMCWRITEDATA(30)",
	OutTemp       => MIMCWRITEDATA_OUT(30),
	Paths         => (0 => (CPMMCCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => MIMCWRITEDATA(31),
	GlitchData    => MIMCWRITEDATA31_GlitchData,
	OutSignalName => "MIMCWRITEDATA(31)",
	OutTemp       => MIMCWRITEDATA_OUT(31),
	Paths         => (0 => (CPMMCCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => MIMCWRITEDATA(32),
	GlitchData    => MIMCWRITEDATA32_GlitchData,
	OutSignalName => "MIMCWRITEDATA(32)",
	OutTemp       => MIMCWRITEDATA_OUT(32),
	Paths         => (0 => (CPMMCCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => MIMCWRITEDATA(33),
	GlitchData    => MIMCWRITEDATA33_GlitchData,
	OutSignalName => "MIMCWRITEDATA(33)",
	OutTemp       => MIMCWRITEDATA_OUT(33),
	Paths         => (0 => (CPMMCCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => MIMCWRITEDATA(34),
	GlitchData    => MIMCWRITEDATA34_GlitchData,
	OutSignalName => "MIMCWRITEDATA(34)",
	OutTemp       => MIMCWRITEDATA_OUT(34),
	Paths         => (0 => (CPMMCCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => MIMCWRITEDATA(35),
	GlitchData    => MIMCWRITEDATA35_GlitchData,
	OutSignalName => "MIMCWRITEDATA(35)",
	OutTemp       => MIMCWRITEDATA_OUT(35),
	Paths         => (0 => (CPMMCCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => MIMCWRITEDATA(36),
	GlitchData    => MIMCWRITEDATA36_GlitchData,
	OutSignalName => "MIMCWRITEDATA(36)",
	OutTemp       => MIMCWRITEDATA_OUT(36),
	Paths         => (0 => (CPMMCCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => MIMCWRITEDATA(37),
	GlitchData    => MIMCWRITEDATA37_GlitchData,
	OutSignalName => "MIMCWRITEDATA(37)",
	OutTemp       => MIMCWRITEDATA_OUT(37),
	Paths         => (0 => (CPMMCCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => MIMCWRITEDATA(38),
	GlitchData    => MIMCWRITEDATA38_GlitchData,
	OutSignalName => "MIMCWRITEDATA(38)",
	OutTemp       => MIMCWRITEDATA_OUT(38),
	Paths         => (0 => (CPMMCCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => MIMCWRITEDATA(39),
	GlitchData    => MIMCWRITEDATA39_GlitchData,
	OutSignalName => "MIMCWRITEDATA(39)",
	OutTemp       => MIMCWRITEDATA_OUT(39),
	Paths         => (0 => (CPMMCCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => MIMCWRITEDATA(40),
	GlitchData    => MIMCWRITEDATA40_GlitchData,
	OutSignalName => "MIMCWRITEDATA(40)",
	OutTemp       => MIMCWRITEDATA_OUT(40),
	Paths         => (0 => (CPMMCCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => MIMCWRITEDATA(41),
	GlitchData    => MIMCWRITEDATA41_GlitchData,
	OutSignalName => "MIMCWRITEDATA(41)",
	OutTemp       => MIMCWRITEDATA_OUT(41),
	Paths         => (0 => (CPMMCCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => MIMCWRITEDATA(42),
	GlitchData    => MIMCWRITEDATA42_GlitchData,
	OutSignalName => "MIMCWRITEDATA(42)",
	OutTemp       => MIMCWRITEDATA_OUT(42),
	Paths         => (0 => (CPMMCCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => MIMCWRITEDATA(43),
	GlitchData    => MIMCWRITEDATA43_GlitchData,
	OutSignalName => "MIMCWRITEDATA(43)",
	OutTemp       => MIMCWRITEDATA_OUT(43),
	Paths         => (0 => (CPMMCCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => MIMCWRITEDATA(44),
	GlitchData    => MIMCWRITEDATA44_GlitchData,
	OutSignalName => "MIMCWRITEDATA(44)",
	OutTemp       => MIMCWRITEDATA_OUT(44),
	Paths         => (0 => (CPMMCCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => MIMCWRITEDATA(45),
	GlitchData    => MIMCWRITEDATA45_GlitchData,
	OutSignalName => "MIMCWRITEDATA(45)",
	OutTemp       => MIMCWRITEDATA_OUT(45),
	Paths         => (0 => (CPMMCCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => MIMCWRITEDATA(46),
	GlitchData    => MIMCWRITEDATA46_GlitchData,
	OutSignalName => "MIMCWRITEDATA(46)",
	OutTemp       => MIMCWRITEDATA_OUT(46),
	Paths         => (0 => (CPMMCCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => MIMCWRITEDATA(47),
	GlitchData    => MIMCWRITEDATA47_GlitchData,
	OutSignalName => "MIMCWRITEDATA(47)",
	OutTemp       => MIMCWRITEDATA_OUT(47),
	Paths         => (0 => (CPMMCCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => MIMCWRITEDATA(48),
	GlitchData    => MIMCWRITEDATA48_GlitchData,
	OutSignalName => "MIMCWRITEDATA(48)",
	OutTemp       => MIMCWRITEDATA_OUT(48),
	Paths         => (0 => (CPMMCCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => MIMCWRITEDATA(49),
	GlitchData    => MIMCWRITEDATA49_GlitchData,
	OutSignalName => "MIMCWRITEDATA(49)",
	OutTemp       => MIMCWRITEDATA_OUT(49),
	Paths         => (0 => (CPMMCCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => MIMCWRITEDATA(50),
	GlitchData    => MIMCWRITEDATA50_GlitchData,
	OutSignalName => "MIMCWRITEDATA(50)",
	OutTemp       => MIMCWRITEDATA_OUT(50),
	Paths         => (0 => (CPMMCCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => MIMCWRITEDATA(51),
	GlitchData    => MIMCWRITEDATA51_GlitchData,
	OutSignalName => "MIMCWRITEDATA(51)",
	OutTemp       => MIMCWRITEDATA_OUT(51),
	Paths         => (0 => (CPMMCCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => MIMCWRITEDATA(52),
	GlitchData    => MIMCWRITEDATA52_GlitchData,
	OutSignalName => "MIMCWRITEDATA(52)",
	OutTemp       => MIMCWRITEDATA_OUT(52),
	Paths         => (0 => (CPMMCCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => MIMCWRITEDATA(53),
	GlitchData    => MIMCWRITEDATA53_GlitchData,
	OutSignalName => "MIMCWRITEDATA(53)",
	OutTemp       => MIMCWRITEDATA_OUT(53),
	Paths         => (0 => (CPMMCCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => MIMCWRITEDATA(54),
	GlitchData    => MIMCWRITEDATA54_GlitchData,
	OutSignalName => "MIMCWRITEDATA(54)",
	OutTemp       => MIMCWRITEDATA_OUT(54),
	Paths         => (0 => (CPMMCCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => MIMCWRITEDATA(55),
	GlitchData    => MIMCWRITEDATA55_GlitchData,
	OutSignalName => "MIMCWRITEDATA(55)",
	OutTemp       => MIMCWRITEDATA_OUT(55),
	Paths         => (0 => (CPMMCCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => MIMCWRITEDATA(56),
	GlitchData    => MIMCWRITEDATA56_GlitchData,
	OutSignalName => "MIMCWRITEDATA(56)",
	OutTemp       => MIMCWRITEDATA_OUT(56),
	Paths         => (0 => (CPMMCCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => MIMCWRITEDATA(57),
	GlitchData    => MIMCWRITEDATA57_GlitchData,
	OutSignalName => "MIMCWRITEDATA(57)",
	OutTemp       => MIMCWRITEDATA_OUT(57),
	Paths         => (0 => (CPMMCCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => MIMCWRITEDATA(58),
	GlitchData    => MIMCWRITEDATA58_GlitchData,
	OutSignalName => "MIMCWRITEDATA(58)",
	OutTemp       => MIMCWRITEDATA_OUT(58),
	Paths         => (0 => (CPMMCCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => MIMCWRITEDATA(59),
	GlitchData    => MIMCWRITEDATA59_GlitchData,
	OutSignalName => "MIMCWRITEDATA(59)",
	OutTemp       => MIMCWRITEDATA_OUT(59),
	Paths         => (0 => (CPMMCCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => MIMCWRITEDATA(60),
	GlitchData    => MIMCWRITEDATA60_GlitchData,
	OutSignalName => "MIMCWRITEDATA(60)",
	OutTemp       => MIMCWRITEDATA_OUT(60),
	Paths         => (0 => (CPMMCCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => MIMCWRITEDATA(61),
	GlitchData    => MIMCWRITEDATA61_GlitchData,
	OutSignalName => "MIMCWRITEDATA(61)",
	OutTemp       => MIMCWRITEDATA_OUT(61),
	Paths         => (0 => (CPMMCCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => MIMCWRITEDATA(62),
	GlitchData    => MIMCWRITEDATA62_GlitchData,
	OutSignalName => "MIMCWRITEDATA(62)",
	OutTemp       => MIMCWRITEDATA_OUT(62),
	Paths         => (0 => (CPMMCCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => MIMCWRITEDATA(63),
	GlitchData    => MIMCWRITEDATA63_GlitchData,
	OutSignalName => "MIMCWRITEDATA(63)",
	OutTemp       => MIMCWRITEDATA_OUT(63),
	Paths         => (0 => (CPMMCCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => MIMCWRITEDATA(64),
	GlitchData    => MIMCWRITEDATA64_GlitchData,
	OutSignalName => "MIMCWRITEDATA(64)",
	OutTemp       => MIMCWRITEDATA_OUT(64),
	Paths         => (0 => (CPMMCCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => MIMCWRITEDATA(65),
	GlitchData    => MIMCWRITEDATA65_GlitchData,
	OutSignalName => "MIMCWRITEDATA(65)",
	OutTemp       => MIMCWRITEDATA_OUT(65),
	Paths         => (0 => (CPMMCCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => MIMCWRITEDATA(66),
	GlitchData    => MIMCWRITEDATA66_GlitchData,
	OutSignalName => "MIMCWRITEDATA(66)",
	OutTemp       => MIMCWRITEDATA_OUT(66),
	Paths         => (0 => (CPMMCCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => MIMCWRITEDATA(67),
	GlitchData    => MIMCWRITEDATA67_GlitchData,
	OutSignalName => "MIMCWRITEDATA(67)",
	OutTemp       => MIMCWRITEDATA_OUT(67),
	Paths         => (0 => (CPMMCCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => MIMCWRITEDATA(68),
	GlitchData    => MIMCWRITEDATA68_GlitchData,
	OutSignalName => "MIMCWRITEDATA(68)",
	OutTemp       => MIMCWRITEDATA_OUT(68),
	Paths         => (0 => (CPMMCCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => MIMCWRITEDATA(69),
	GlitchData    => MIMCWRITEDATA69_GlitchData,
	OutSignalName => "MIMCWRITEDATA(69)",
	OutTemp       => MIMCWRITEDATA_OUT(69),
	Paths         => (0 => (CPMMCCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => MIMCWRITEDATA(70),
	GlitchData    => MIMCWRITEDATA70_GlitchData,
	OutSignalName => "MIMCWRITEDATA(70)",
	OutTemp       => MIMCWRITEDATA_OUT(70),
	Paths         => (0 => (CPMMCCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => MIMCWRITEDATA(71),
	GlitchData    => MIMCWRITEDATA71_GlitchData,
	OutSignalName => "MIMCWRITEDATA(71)",
	OutTemp       => MIMCWRITEDATA_OUT(71),
	Paths         => (0 => (CPMMCCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => MIMCWRITEDATA(72),
	GlitchData    => MIMCWRITEDATA72_GlitchData,
	OutSignalName => "MIMCWRITEDATA(72)",
	OutTemp       => MIMCWRITEDATA_OUT(72),
	Paths         => (0 => (CPMMCCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => MIMCWRITEDATA(73),
	GlitchData    => MIMCWRITEDATA73_GlitchData,
	OutSignalName => "MIMCWRITEDATA(73)",
	OutTemp       => MIMCWRITEDATA_OUT(73),
	Paths         => (0 => (CPMMCCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => MIMCWRITEDATA(74),
	GlitchData    => MIMCWRITEDATA74_GlitchData,
	OutSignalName => "MIMCWRITEDATA(74)",
	OutTemp       => MIMCWRITEDATA_OUT(74),
	Paths         => (0 => (CPMMCCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => MIMCWRITEDATA(75),
	GlitchData    => MIMCWRITEDATA75_GlitchData,
	OutSignalName => "MIMCWRITEDATA(75)",
	OutTemp       => MIMCWRITEDATA_OUT(75),
	Paths         => (0 => (CPMMCCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => MIMCWRITEDATA(76),
	GlitchData    => MIMCWRITEDATA76_GlitchData,
	OutSignalName => "MIMCWRITEDATA(76)",
	OutTemp       => MIMCWRITEDATA_OUT(76),
	Paths         => (0 => (CPMMCCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => MIMCWRITEDATA(77),
	GlitchData    => MIMCWRITEDATA77_GlitchData,
	OutSignalName => "MIMCWRITEDATA(77)",
	OutTemp       => MIMCWRITEDATA_OUT(77),
	Paths         => (0 => (CPMMCCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => MIMCWRITEDATA(78),
	GlitchData    => MIMCWRITEDATA78_GlitchData,
	OutSignalName => "MIMCWRITEDATA(78)",
	OutTemp       => MIMCWRITEDATA_OUT(78),
	Paths         => (0 => (CPMMCCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => MIMCWRITEDATA(79),
	GlitchData    => MIMCWRITEDATA79_GlitchData,
	OutSignalName => "MIMCWRITEDATA(79)",
	OutTemp       => MIMCWRITEDATA_OUT(79),
	Paths         => (0 => (CPMMCCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => MIMCWRITEDATA(80),
	GlitchData    => MIMCWRITEDATA80_GlitchData,
	OutSignalName => "MIMCWRITEDATA(80)",
	OutTemp       => MIMCWRITEDATA_OUT(80),
	Paths         => (0 => (CPMMCCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => MIMCWRITEDATA(81),
	GlitchData    => MIMCWRITEDATA81_GlitchData,
	OutSignalName => "MIMCWRITEDATA(81)",
	OutTemp       => MIMCWRITEDATA_OUT(81),
	Paths         => (0 => (CPMMCCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => MIMCWRITEDATA(82),
	GlitchData    => MIMCWRITEDATA82_GlitchData,
	OutSignalName => "MIMCWRITEDATA(82)",
	OutTemp       => MIMCWRITEDATA_OUT(82),
	Paths         => (0 => (CPMMCCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => MIMCWRITEDATA(83),
	GlitchData    => MIMCWRITEDATA83_GlitchData,
	OutSignalName => "MIMCWRITEDATA(83)",
	OutTemp       => MIMCWRITEDATA_OUT(83),
	Paths         => (0 => (CPMMCCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => MIMCWRITEDATA(84),
	GlitchData    => MIMCWRITEDATA84_GlitchData,
	OutSignalName => "MIMCWRITEDATA(84)",
	OutTemp       => MIMCWRITEDATA_OUT(84),
	Paths         => (0 => (CPMMCCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => MIMCWRITEDATA(85),
	GlitchData    => MIMCWRITEDATA85_GlitchData,
	OutSignalName => "MIMCWRITEDATA(85)",
	OutTemp       => MIMCWRITEDATA_OUT(85),
	Paths         => (0 => (CPMMCCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => MIMCWRITEDATA(86),
	GlitchData    => MIMCWRITEDATA86_GlitchData,
	OutSignalName => "MIMCWRITEDATA(86)",
	OutTemp       => MIMCWRITEDATA_OUT(86),
	Paths         => (0 => (CPMMCCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => MIMCWRITEDATA(87),
	GlitchData    => MIMCWRITEDATA87_GlitchData,
	OutSignalName => "MIMCWRITEDATA(87)",
	OutTemp       => MIMCWRITEDATA_OUT(87),
	Paths         => (0 => (CPMMCCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => MIMCWRITEDATA(88),
	GlitchData    => MIMCWRITEDATA88_GlitchData,
	OutSignalName => "MIMCWRITEDATA(88)",
	OutTemp       => MIMCWRITEDATA_OUT(88),
	Paths         => (0 => (CPMMCCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => MIMCWRITEDATA(89),
	GlitchData    => MIMCWRITEDATA89_GlitchData,
	OutSignalName => "MIMCWRITEDATA(89)",
	OutTemp       => MIMCWRITEDATA_OUT(89),
	Paths         => (0 => (CPMMCCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => MIMCWRITEDATA(90),
	GlitchData    => MIMCWRITEDATA90_GlitchData,
	OutSignalName => "MIMCWRITEDATA(90)",
	OutTemp       => MIMCWRITEDATA_OUT(90),
	Paths         => (0 => (CPMMCCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => MIMCWRITEDATA(91),
	GlitchData    => MIMCWRITEDATA91_GlitchData,
	OutSignalName => "MIMCWRITEDATA(91)",
	OutTemp       => MIMCWRITEDATA_OUT(91),
	Paths         => (0 => (CPMMCCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => MIMCWRITEDATA(92),
	GlitchData    => MIMCWRITEDATA92_GlitchData,
	OutSignalName => "MIMCWRITEDATA(92)",
	OutTemp       => MIMCWRITEDATA_OUT(92),
	Paths         => (0 => (CPMMCCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => MIMCWRITEDATA(93),
	GlitchData    => MIMCWRITEDATA93_GlitchData,
	OutSignalName => "MIMCWRITEDATA(93)",
	OutTemp       => MIMCWRITEDATA_OUT(93),
	Paths         => (0 => (CPMMCCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => MIMCWRITEDATA(94),
	GlitchData    => MIMCWRITEDATA94_GlitchData,
	OutSignalName => "MIMCWRITEDATA(94)",
	OutTemp       => MIMCWRITEDATA_OUT(94),
	Paths         => (0 => (CPMMCCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => MIMCWRITEDATA(95),
	GlitchData    => MIMCWRITEDATA95_GlitchData,
	OutSignalName => "MIMCWRITEDATA(95)",
	OutTemp       => MIMCWRITEDATA_OUT(95),
	Paths         => (0 => (CPMMCCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => MIMCWRITEDATA(96),
	GlitchData    => MIMCWRITEDATA96_GlitchData,
	OutSignalName => "MIMCWRITEDATA(96)",
	OutTemp       => MIMCWRITEDATA_OUT(96),
	Paths         => (0 => (CPMMCCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => MIMCWRITEDATA(97),
	GlitchData    => MIMCWRITEDATA97_GlitchData,
	OutSignalName => "MIMCWRITEDATA(97)",
	OutTemp       => MIMCWRITEDATA_OUT(97),
	Paths         => (0 => (CPMMCCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => MIMCWRITEDATA(98),
	GlitchData    => MIMCWRITEDATA98_GlitchData,
	OutSignalName => "MIMCWRITEDATA(98)",
	OutTemp       => MIMCWRITEDATA_OUT(98),
	Paths         => (0 => (CPMMCCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => MIMCWRITEDATA(99),
	GlitchData    => MIMCWRITEDATA99_GlitchData,
	OutSignalName => "MIMCWRITEDATA(99)",
	OutTemp       => MIMCWRITEDATA_OUT(99),
	Paths         => (0 => (CPMMCCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => MIMCWRITEDATA(100),
	GlitchData    => MIMCWRITEDATA100_GlitchData,
	OutSignalName => "MIMCWRITEDATA(100)",
	OutTemp       => MIMCWRITEDATA_OUT(100),
	Paths         => (0 => (CPMMCCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => MIMCWRITEDATA(101),
	GlitchData    => MIMCWRITEDATA101_GlitchData,
	OutSignalName => "MIMCWRITEDATA(101)",
	OutTemp       => MIMCWRITEDATA_OUT(101),
	Paths         => (0 => (CPMMCCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => MIMCWRITEDATA(102),
	GlitchData    => MIMCWRITEDATA102_GlitchData,
	OutSignalName => "MIMCWRITEDATA(102)",
	OutTemp       => MIMCWRITEDATA_OUT(102),
	Paths         => (0 => (CPMMCCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => MIMCWRITEDATA(103),
	GlitchData    => MIMCWRITEDATA103_GlitchData,
	OutSignalName => "MIMCWRITEDATA(103)",
	OutTemp       => MIMCWRITEDATA_OUT(103),
	Paths         => (0 => (CPMMCCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => MIMCWRITEDATA(104),
	GlitchData    => MIMCWRITEDATA104_GlitchData,
	OutSignalName => "MIMCWRITEDATA(104)",
	OutTemp       => MIMCWRITEDATA_OUT(104),
	Paths         => (0 => (CPMMCCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => MIMCWRITEDATA(105),
	GlitchData    => MIMCWRITEDATA105_GlitchData,
	OutSignalName => "MIMCWRITEDATA(105)",
	OutTemp       => MIMCWRITEDATA_OUT(105),
	Paths         => (0 => (CPMMCCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => MIMCWRITEDATA(106),
	GlitchData    => MIMCWRITEDATA106_GlitchData,
	OutSignalName => "MIMCWRITEDATA(106)",
	OutTemp       => MIMCWRITEDATA_OUT(106),
	Paths         => (0 => (CPMMCCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => MIMCWRITEDATA(107),
	GlitchData    => MIMCWRITEDATA107_GlitchData,
	OutSignalName => "MIMCWRITEDATA(107)",
	OutTemp       => MIMCWRITEDATA_OUT(107),
	Paths         => (0 => (CPMMCCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => MIMCWRITEDATA(108),
	GlitchData    => MIMCWRITEDATA108_GlitchData,
	OutSignalName => "MIMCWRITEDATA(108)",
	OutTemp       => MIMCWRITEDATA_OUT(108),
	Paths         => (0 => (CPMMCCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => MIMCWRITEDATA(109),
	GlitchData    => MIMCWRITEDATA109_GlitchData,
	OutSignalName => "MIMCWRITEDATA(109)",
	OutTemp       => MIMCWRITEDATA_OUT(109),
	Paths         => (0 => (CPMMCCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => MIMCWRITEDATA(110),
	GlitchData    => MIMCWRITEDATA110_GlitchData,
	OutSignalName => "MIMCWRITEDATA(110)",
	OutTemp       => MIMCWRITEDATA_OUT(110),
	Paths         => (0 => (CPMMCCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => MIMCWRITEDATA(111),
	GlitchData    => MIMCWRITEDATA111_GlitchData,
	OutSignalName => "MIMCWRITEDATA(111)",
	OutTemp       => MIMCWRITEDATA_OUT(111),
	Paths         => (0 => (CPMMCCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => MIMCWRITEDATA(112),
	GlitchData    => MIMCWRITEDATA112_GlitchData,
	OutSignalName => "MIMCWRITEDATA(112)",
	OutTemp       => MIMCWRITEDATA_OUT(112),
	Paths         => (0 => (CPMMCCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => MIMCWRITEDATA(113),
	GlitchData    => MIMCWRITEDATA113_GlitchData,
	OutSignalName => "MIMCWRITEDATA(113)",
	OutTemp       => MIMCWRITEDATA_OUT(113),
	Paths         => (0 => (CPMMCCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => MIMCWRITEDATA(114),
	GlitchData    => MIMCWRITEDATA114_GlitchData,
	OutSignalName => "MIMCWRITEDATA(114)",
	OutTemp       => MIMCWRITEDATA_OUT(114),
	Paths         => (0 => (CPMMCCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => MIMCWRITEDATA(115),
	GlitchData    => MIMCWRITEDATA115_GlitchData,
	OutSignalName => "MIMCWRITEDATA(115)",
	OutTemp       => MIMCWRITEDATA_OUT(115),
	Paths         => (0 => (CPMMCCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => MIMCWRITEDATA(116),
	GlitchData    => MIMCWRITEDATA116_GlitchData,
	OutSignalName => "MIMCWRITEDATA(116)",
	OutTemp       => MIMCWRITEDATA_OUT(116),
	Paths         => (0 => (CPMMCCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => MIMCWRITEDATA(117),
	GlitchData    => MIMCWRITEDATA117_GlitchData,
	OutSignalName => "MIMCWRITEDATA(117)",
	OutTemp       => MIMCWRITEDATA_OUT(117),
	Paths         => (0 => (CPMMCCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => MIMCWRITEDATA(118),
	GlitchData    => MIMCWRITEDATA118_GlitchData,
	OutSignalName => "MIMCWRITEDATA(118)",
	OutTemp       => MIMCWRITEDATA_OUT(118),
	Paths         => (0 => (CPMMCCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => MIMCWRITEDATA(119),
	GlitchData    => MIMCWRITEDATA119_GlitchData,
	OutSignalName => "MIMCWRITEDATA(119)",
	OutTemp       => MIMCWRITEDATA_OUT(119),
	Paths         => (0 => (CPMMCCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => MIMCWRITEDATA(120),
	GlitchData    => MIMCWRITEDATA120_GlitchData,
	OutSignalName => "MIMCWRITEDATA(120)",
	OutTemp       => MIMCWRITEDATA_OUT(120),
	Paths         => (0 => (CPMMCCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => MIMCWRITEDATA(121),
	GlitchData    => MIMCWRITEDATA121_GlitchData,
	OutSignalName => "MIMCWRITEDATA(121)",
	OutTemp       => MIMCWRITEDATA_OUT(121),
	Paths         => (0 => (CPMMCCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => MIMCWRITEDATA(122),
	GlitchData    => MIMCWRITEDATA122_GlitchData,
	OutSignalName => "MIMCWRITEDATA(122)",
	OutTemp       => MIMCWRITEDATA_OUT(122),
	Paths         => (0 => (CPMMCCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => MIMCWRITEDATA(123),
	GlitchData    => MIMCWRITEDATA123_GlitchData,
	OutSignalName => "MIMCWRITEDATA(123)",
	OutTemp       => MIMCWRITEDATA_OUT(123),
	Paths         => (0 => (CPMMCCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => MIMCWRITEDATA(124),
	GlitchData    => MIMCWRITEDATA124_GlitchData,
	OutSignalName => "MIMCWRITEDATA(124)",
	OutTemp       => MIMCWRITEDATA_OUT(124),
	Paths         => (0 => (CPMMCCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => MIMCWRITEDATA(125),
	GlitchData    => MIMCWRITEDATA125_GlitchData,
	OutSignalName => "MIMCWRITEDATA(125)",
	OutTemp       => MIMCWRITEDATA_OUT(125),
	Paths         => (0 => (CPMMCCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => MIMCWRITEDATA(126),
	GlitchData    => MIMCWRITEDATA126_GlitchData,
	OutSignalName => "MIMCWRITEDATA(126)",
	OutTemp       => MIMCWRITEDATA_OUT(126),
	Paths         => (0 => (CPMMCCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => MIMCWRITEDATA(127),
	GlitchData    => MIMCWRITEDATA127_GlitchData,
	OutSignalName => "MIMCWRITEDATA(127)",
	OutTemp       => MIMCWRITEDATA_OUT(127),
	Paths         => (0 => (CPMMCCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => MIMCWRITEDATAVALID,
	GlitchData    => MIMCWRITEDATAVALID_GlitchData,
	OutSignalName => "MIMCWRITEDATAVALID",
	OutTemp       => MIMCWRITEDATAVALID_OUT,
	Paths         => (0 => (CPMMCCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCCPMINTERCONNECTBUSY,
	GlitchData    => PPCCPMINTERCONNECTBUSY_GlitchData,
	OutSignalName => "PPCCPMINTERCONNECTBUSY",
	OutTemp       => PPCCPMINTERCONNECTBUSY_OUT,
	Paths         => (0 => (CPMINTERCONNECTCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCDSDCRACK,
	GlitchData    => PPCDSDCRACK_GlitchData,
	OutSignalName => "PPCDSDCRACK",
	OutTemp       => PPCDSDCRACK_OUT,
	Paths         => (0 => (CPMDCRCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCDSDCRTIMEOUTWAIT,
	GlitchData    => PPCDSDCRTIMEOUTWAIT_GlitchData,
	OutSignalName => "PPCDSDCRTIMEOUTWAIT",
	OutTemp       => PPCDSDCRTIMEOUTWAIT_OUT,
	Paths         => (0 => (CPMDCRCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCDSDCRDBUSIN(0),
	GlitchData    => PPCDSDCRDBUSIN0_GlitchData,
	OutSignalName => "PPCDSDCRDBUSIN(0)",
	OutTemp       => PPCDSDCRDBUSIN_OUT(0),
	Paths         => (0 => (CPMDCRCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCDSDCRDBUSIN(1),
	GlitchData    => PPCDSDCRDBUSIN1_GlitchData,
	OutSignalName => "PPCDSDCRDBUSIN(1)",
	OutTemp       => PPCDSDCRDBUSIN_OUT(1),
	Paths         => (0 => (CPMDCRCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCDSDCRDBUSIN(2),
	GlitchData    => PPCDSDCRDBUSIN2_GlitchData,
	OutSignalName => "PPCDSDCRDBUSIN(2)",
	OutTemp       => PPCDSDCRDBUSIN_OUT(2),
	Paths         => (0 => (CPMDCRCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCDSDCRDBUSIN(3),
	GlitchData    => PPCDSDCRDBUSIN3_GlitchData,
	OutSignalName => "PPCDSDCRDBUSIN(3)",
	OutTemp       => PPCDSDCRDBUSIN_OUT(3),
	Paths         => (0 => (CPMDCRCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCDSDCRDBUSIN(4),
	GlitchData    => PPCDSDCRDBUSIN4_GlitchData,
	OutSignalName => "PPCDSDCRDBUSIN(4)",
	OutTemp       => PPCDSDCRDBUSIN_OUT(4),
	Paths         => (0 => (CPMDCRCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCDSDCRDBUSIN(5),
	GlitchData    => PPCDSDCRDBUSIN5_GlitchData,
	OutSignalName => "PPCDSDCRDBUSIN(5)",
	OutTemp       => PPCDSDCRDBUSIN_OUT(5),
	Paths         => (0 => (CPMDCRCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCDSDCRDBUSIN(6),
	GlitchData    => PPCDSDCRDBUSIN6_GlitchData,
	OutSignalName => "PPCDSDCRDBUSIN(6)",
	OutTemp       => PPCDSDCRDBUSIN_OUT(6),
	Paths         => (0 => (CPMDCRCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCDSDCRDBUSIN(7),
	GlitchData    => PPCDSDCRDBUSIN7_GlitchData,
	OutSignalName => "PPCDSDCRDBUSIN(7)",
	OutTemp       => PPCDSDCRDBUSIN_OUT(7),
	Paths         => (0 => (CPMDCRCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCDSDCRDBUSIN(8),
	GlitchData    => PPCDSDCRDBUSIN8_GlitchData,
	OutSignalName => "PPCDSDCRDBUSIN(8)",
	OutTemp       => PPCDSDCRDBUSIN_OUT(8),
	Paths         => (0 => (CPMDCRCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCDSDCRDBUSIN(9),
	GlitchData    => PPCDSDCRDBUSIN9_GlitchData,
	OutSignalName => "PPCDSDCRDBUSIN(9)",
	OutTemp       => PPCDSDCRDBUSIN_OUT(9),
	Paths         => (0 => (CPMDCRCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCDSDCRDBUSIN(10),
	GlitchData    => PPCDSDCRDBUSIN10_GlitchData,
	OutSignalName => "PPCDSDCRDBUSIN(10)",
	OutTemp       => PPCDSDCRDBUSIN_OUT(10),
	Paths         => (0 => (CPMDCRCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCDSDCRDBUSIN(11),
	GlitchData    => PPCDSDCRDBUSIN11_GlitchData,
	OutSignalName => "PPCDSDCRDBUSIN(11)",
	OutTemp       => PPCDSDCRDBUSIN_OUT(11),
	Paths         => (0 => (CPMDCRCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCDSDCRDBUSIN(12),
	GlitchData    => PPCDSDCRDBUSIN12_GlitchData,
	OutSignalName => "PPCDSDCRDBUSIN(12)",
	OutTemp       => PPCDSDCRDBUSIN_OUT(12),
	Paths         => (0 => (CPMDCRCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCDSDCRDBUSIN(13),
	GlitchData    => PPCDSDCRDBUSIN13_GlitchData,
	OutSignalName => "PPCDSDCRDBUSIN(13)",
	OutTemp       => PPCDSDCRDBUSIN_OUT(13),
	Paths         => (0 => (CPMDCRCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCDSDCRDBUSIN(14),
	GlitchData    => PPCDSDCRDBUSIN14_GlitchData,
	OutSignalName => "PPCDSDCRDBUSIN(14)",
	OutTemp       => PPCDSDCRDBUSIN_OUT(14),
	Paths         => (0 => (CPMDCRCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCDSDCRDBUSIN(15),
	GlitchData    => PPCDSDCRDBUSIN15_GlitchData,
	OutSignalName => "PPCDSDCRDBUSIN(15)",
	OutTemp       => PPCDSDCRDBUSIN_OUT(15),
	Paths         => (0 => (CPMDCRCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCDSDCRDBUSIN(16),
	GlitchData    => PPCDSDCRDBUSIN16_GlitchData,
	OutSignalName => "PPCDSDCRDBUSIN(16)",
	OutTemp       => PPCDSDCRDBUSIN_OUT(16),
	Paths         => (0 => (CPMDCRCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCDSDCRDBUSIN(17),
	GlitchData    => PPCDSDCRDBUSIN17_GlitchData,
	OutSignalName => "PPCDSDCRDBUSIN(17)",
	OutTemp       => PPCDSDCRDBUSIN_OUT(17),
	Paths         => (0 => (CPMDCRCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCDSDCRDBUSIN(18),
	GlitchData    => PPCDSDCRDBUSIN18_GlitchData,
	OutSignalName => "PPCDSDCRDBUSIN(18)",
	OutTemp       => PPCDSDCRDBUSIN_OUT(18),
	Paths         => (0 => (CPMDCRCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCDSDCRDBUSIN(19),
	GlitchData    => PPCDSDCRDBUSIN19_GlitchData,
	OutSignalName => "PPCDSDCRDBUSIN(19)",
	OutTemp       => PPCDSDCRDBUSIN_OUT(19),
	Paths         => (0 => (CPMDCRCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCDSDCRDBUSIN(20),
	GlitchData    => PPCDSDCRDBUSIN20_GlitchData,
	OutSignalName => "PPCDSDCRDBUSIN(20)",
	OutTemp       => PPCDSDCRDBUSIN_OUT(20),
	Paths         => (0 => (CPMDCRCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCDSDCRDBUSIN(21),
	GlitchData    => PPCDSDCRDBUSIN21_GlitchData,
	OutSignalName => "PPCDSDCRDBUSIN(21)",
	OutTemp       => PPCDSDCRDBUSIN_OUT(21),
	Paths         => (0 => (CPMDCRCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCDSDCRDBUSIN(22),
	GlitchData    => PPCDSDCRDBUSIN22_GlitchData,
	OutSignalName => "PPCDSDCRDBUSIN(22)",
	OutTemp       => PPCDSDCRDBUSIN_OUT(22),
	Paths         => (0 => (CPMDCRCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCDSDCRDBUSIN(23),
	GlitchData    => PPCDSDCRDBUSIN23_GlitchData,
	OutSignalName => "PPCDSDCRDBUSIN(23)",
	OutTemp       => PPCDSDCRDBUSIN_OUT(23),
	Paths         => (0 => (CPMDCRCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCDSDCRDBUSIN(24),
	GlitchData    => PPCDSDCRDBUSIN24_GlitchData,
	OutSignalName => "PPCDSDCRDBUSIN(24)",
	OutTemp       => PPCDSDCRDBUSIN_OUT(24),
	Paths         => (0 => (CPMDCRCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCDSDCRDBUSIN(25),
	GlitchData    => PPCDSDCRDBUSIN25_GlitchData,
	OutSignalName => "PPCDSDCRDBUSIN(25)",
	OutTemp       => PPCDSDCRDBUSIN_OUT(25),
	Paths         => (0 => (CPMDCRCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCDSDCRDBUSIN(26),
	GlitchData    => PPCDSDCRDBUSIN26_GlitchData,
	OutSignalName => "PPCDSDCRDBUSIN(26)",
	OutTemp       => PPCDSDCRDBUSIN_OUT(26),
	Paths         => (0 => (CPMDCRCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCDSDCRDBUSIN(27),
	GlitchData    => PPCDSDCRDBUSIN27_GlitchData,
	OutSignalName => "PPCDSDCRDBUSIN(27)",
	OutTemp       => PPCDSDCRDBUSIN_OUT(27),
	Paths         => (0 => (CPMDCRCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCDSDCRDBUSIN(28),
	GlitchData    => PPCDSDCRDBUSIN28_GlitchData,
	OutSignalName => "PPCDSDCRDBUSIN(28)",
	OutTemp       => PPCDSDCRDBUSIN_OUT(28),
	Paths         => (0 => (CPMDCRCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCDSDCRDBUSIN(29),
	GlitchData    => PPCDSDCRDBUSIN29_GlitchData,
	OutSignalName => "PPCDSDCRDBUSIN(29)",
	OutTemp       => PPCDSDCRDBUSIN_OUT(29),
	Paths         => (0 => (CPMDCRCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCDSDCRDBUSIN(30),
	GlitchData    => PPCDSDCRDBUSIN30_GlitchData,
	OutSignalName => "PPCDSDCRDBUSIN(30)",
	OutTemp       => PPCDSDCRDBUSIN_OUT(30),
	Paths         => (0 => (CPMDCRCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCDSDCRDBUSIN(31),
	GlitchData    => PPCDSDCRDBUSIN31_GlitchData,
	OutSignalName => "PPCDSDCRDBUSIN(31)",
	OutTemp       => PPCDSDCRDBUSIN_OUT(31),
	Paths         => (0 => (CPMDCRCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCEICINTERCONNECTIRQ,
	GlitchData    => PPCEICINTERCONNECTIRQ_GlitchData,
	OutSignalName => "PPCEICINTERCONNECTIRQ",
	OutTemp       => PPCEICINTERCONNECTIRQ_OUT,
	Paths         => (0 => (CPMINTERCONNECTCLK_ipd'last_event, PATH_DELAY,TRUE)),
	Mode          => VitalTransport, DefaultDelay  => PATH_DELAY,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);

   wait on
	APUFCMDECFPUOP_out,
	APUFCMDECLDSTXFERSIZE_out,
	APUFCMDECLOAD_out,
	APUFCMDECNONAUTON_out,
	APUFCMDECSTORE_out,
	APUFCMDECUDIVALID_out,
	APUFCMDECUDI_out,
	APUFCMENDIAN_out,
	APUFCMFLUSH_out,
	APUFCMINSTRUCTION_out,
	APUFCMINSTRVALID_out,
	APUFCMLOADBYTEADDR_out,
	APUFCMLOADDATA_out,
	APUFCMLOADDVALID_out,
	APUFCMMSRFE0_out,
	APUFCMMSRFE1_out,
	APUFCMNEXTINSTRREADY_out,
	APUFCMOPERANDVALID_out,
	APUFCMRADATA_out,
	APUFCMRBDATA_out,
	APUFCMWRITEBACKOK_out,
	C440CPMCORESLEEPREQ_out,
	C440CPMDECIRPTREQ_out,
	C440CPMFITIRPTREQ_out,
	C440CPMMSRCE_out,
	C440CPMMSREE_out,
	C440CPMTIMERRESETREQ_out,
	C440CPMWDIRPTREQ_out,
	C440DBGSYSTEMCONTROL_out,
	C440JTGTDOEN_out,
	C440JTGTDO_out,
	C440MACHINECHECK_out,
	C440RSTCHIPRESETREQ_out,
	C440RSTCORERESETREQ_out,
	C440RSTSYSTEMRESETREQ_out,
	C440TRCBRANCHSTATUS_out,
	C440TRCCYCLE_out,
	C440TRCEXECUTIONSTATUS_out,
	C440TRCTRACESTATUS_out,
	C440TRCTRIGGEREVENTOUT_out,
	C440TRCTRIGGEREVENTTYPE_out,
	DMA0LLRSTENGINEACK_out,
	DMA0LLRXDSTRDYN_out,
	DMA0LLTXD_out,
	DMA0LLTXEOFN_out,
	DMA0LLTXEOPN_out,
	DMA0LLTXREM_out,
	DMA0LLTXSOFN_out,
	DMA0LLTXSOPN_out,
	DMA0LLTXSRCRDYN_out,
	DMA0RXIRQ_out,
	DMA0TXIRQ_out,
	DMA1LLRSTENGINEACK_out,
	DMA1LLRXDSTRDYN_out,
	DMA1LLTXD_out,
	DMA1LLTXEOFN_out,
	DMA1LLTXEOPN_out,
	DMA1LLTXREM_out,
	DMA1LLTXSOFN_out,
	DMA1LLTXSOPN_out,
	DMA1LLTXSRCRDYN_out,
	DMA1RXIRQ_out,
	DMA1TXIRQ_out,
	DMA2LLRSTENGINEACK_out,
	DMA2LLRXDSTRDYN_out,
	DMA2LLTXD_out,
	DMA2LLTXEOFN_out,
	DMA2LLTXEOPN_out,
	DMA2LLTXREM_out,
	DMA2LLTXSOFN_out,
	DMA2LLTXSOPN_out,
	DMA2LLTXSRCRDYN_out,
	DMA2RXIRQ_out,
	DMA2TXIRQ_out,
	DMA3LLRSTENGINEACK_out,
	DMA3LLRXDSTRDYN_out,
	DMA3LLTXD_out,
	DMA3LLTXEOFN_out,
	DMA3LLTXEOPN_out,
	DMA3LLTXREM_out,
	DMA3LLTXSOFN_out,
	DMA3LLTXSOPN_out,
	DMA3LLTXSRCRDYN_out,
	DMA3RXIRQ_out,
	DMA3TXIRQ_out,
	MIMCADDRESSVALID_out,
	MIMCADDRESS_out,
	MIMCBANKCONFLICT_out,
	MIMCBYTEENABLE_out,
	MIMCREADNOTWRITE_out,
	MIMCROWCONFLICT_out,
	MIMCWRITEDATAVALID_out,
	MIMCWRITEDATA_out,
	PPCCPMINTERCONNECTBUSY_out,
	PPCDMDCRABUS_out,
	PPCDMDCRDBUSOUT_out,
	PPCDMDCRREAD_out,
	PPCDMDCRUABUS_out,
	PPCDMDCRWRITE_out,
	PPCDSDCRACK_out,
	PPCDSDCRDBUSIN_out,
	PPCDSDCRTIMEOUTWAIT_out,
	PPCEICINTERCONNECTIRQ_out,
	PPCMPLBABORT_out,
	PPCMPLBABUS_out,
	PPCMPLBBE_out,
	PPCMPLBBUSLOCK_out,
	PPCMPLBLOCKERR_out,
	PPCMPLBPRIORITY_out,
	PPCMPLBRDBURST_out,
	PPCMPLBREQUEST_out,
	PPCMPLBRNW_out,
	PPCMPLBSIZE_out,
	PPCMPLBTATTRIBUTE_out,
	PPCMPLBTYPE_out,
	PPCMPLBUABUS_out,
	PPCMPLBWRBURST_out,
	PPCMPLBWRDBUS_out,
	PPCS0PLBADDRACK_out,
	PPCS0PLBMBUSY_out,
	PPCS0PLBMIRQ_out,
	PPCS0PLBMRDERR_out,
	PPCS0PLBMWRERR_out,
	PPCS0PLBRDBTERM_out,
	PPCS0PLBRDCOMP_out,
	PPCS0PLBRDDACK_out,
	PPCS0PLBRDDBUS_out,
	PPCS0PLBRDWDADDR_out,
	PPCS0PLBREARBITRATE_out,
	PPCS0PLBSSIZE_out,
	PPCS0PLBWAIT_out,
	PPCS0PLBWRBTERM_out,
	PPCS0PLBWRCOMP_out,
	PPCS0PLBWRDACK_out,
	PPCS1PLBADDRACK_out,
	PPCS1PLBMBUSY_out,
	PPCS1PLBMIRQ_out,
	PPCS1PLBMRDERR_out,
	PPCS1PLBMWRERR_out,
	PPCS1PLBRDBTERM_out,
	PPCS1PLBRDCOMP_out,
	PPCS1PLBRDDACK_out,
	PPCS1PLBRDDBUS_out,
	PPCS1PLBRDWDADDR_out,
	PPCS1PLBREARBITRATE_out,
	PPCS1PLBSSIZE_out,
	PPCS1PLBWAIT_out,
	PPCS1PLBWRBTERM_out,
	PPCS1PLBWRCOMP_out,
	PPCS1PLBWRDACK_out,

	CPMC440CLKEN_ipd,
	CPMC440CLK_ipd,
	CPMC440CORECLOCKINACTIVE_ipd,
	CPMC440TIMERCLOCK_ipd,
	CPMDCRCLK_ipd,
	CPMDMA0LLCLK_ipd,
	CPMDMA1LLCLK_ipd,
	CPMDMA2LLCLK_ipd,
	CPMDMA3LLCLK_ipd,
	CPMFCMCLK_ipd,
	CPMINTERCONNECTCLKEN_ipd,
	CPMINTERCONNECTCLKNTO1_ipd,
	CPMINTERCONNECTCLK_ipd,
	CPMMCCLK_ipd,
	CPMPPCMPLBCLK_ipd,
	CPMPPCS0PLBCLK_ipd,
	CPMPPCS1PLBCLK_ipd,
	DBGC440DEBUGHALT_ipd,
	DBGC440SYSTEMSTATUS_ipd,
	DBGC440UNCONDDEBUGEVENT_ipd,
	DCRPPCDMACK_ipd,
	DCRPPCDMDBUSIN_ipd,
	DCRPPCDMTIMEOUTWAIT_ipd,
	DCRPPCDSABUS_ipd,
	DCRPPCDSDBUSOUT_ipd,
	DCRPPCDSREAD_ipd,
	DCRPPCDSWRITE_ipd,
	EICC440CRITIRQ_ipd,
	EICC440EXTIRQ_ipd,
	FCMAPUCONFIRMINSTR_ipd,
	FCMAPUCR_ipd,
	FCMAPUDONE_ipd,
	FCMAPUEXCEPTION_ipd,
	FCMAPUFPSCRFEX_ipd,
	FCMAPURESULTVALID_ipd,
	FCMAPURESULT_ipd,
	FCMAPUSLEEPNOTREADY_ipd,
	FCMAPUSTOREDATA_ipd,
	JTGC440TCK_ipd,
	JTGC440TDI_ipd,
	JTGC440TMS_ipd,
	JTGC440TRSTNEG_ipd,
	LLDMA0RSTENGINEREQ_ipd,
	LLDMA0RXD_ipd,
	LLDMA0RXEOFN_ipd,
	LLDMA0RXEOPN_ipd,
	LLDMA0RXREM_ipd,
	LLDMA0RXSOFN_ipd,
	LLDMA0RXSOPN_ipd,
	LLDMA0RXSRCRDYN_ipd,
	LLDMA0TXDSTRDYN_ipd,
	LLDMA1RSTENGINEREQ_ipd,
	LLDMA1RXD_ipd,
	LLDMA1RXEOFN_ipd,
	LLDMA1RXEOPN_ipd,
	LLDMA1RXREM_ipd,
	LLDMA1RXSOFN_ipd,
	LLDMA1RXSOPN_ipd,
	LLDMA1RXSRCRDYN_ipd,
	LLDMA1TXDSTRDYN_ipd,
	LLDMA2RSTENGINEREQ_ipd,
	LLDMA2RXD_ipd,
	LLDMA2RXEOFN_ipd,
	LLDMA2RXEOPN_ipd,
	LLDMA2RXREM_ipd,
	LLDMA2RXSOFN_ipd,
	LLDMA2RXSOPN_ipd,
	LLDMA2RXSRCRDYN_ipd,
	LLDMA2TXDSTRDYN_ipd,
	LLDMA3RSTENGINEREQ_ipd,
	LLDMA3RXD_ipd,
	LLDMA3RXEOFN_ipd,
	LLDMA3RXEOPN_ipd,
	LLDMA3RXREM_ipd,
	LLDMA3RXSOFN_ipd,
	LLDMA3RXSOPN_ipd,
	LLDMA3RXSRCRDYN_ipd,
	LLDMA3TXDSTRDYN_ipd,
	MCMIADDRREADYTOACCEPT_ipd,
	MCMIREADDATAERR_ipd,
	MCMIREADDATAVALID_ipd,
	MCMIREADDATA_ipd,
	PLBPPCMADDRACK_ipd,
	PLBPPCMMBUSY_ipd,
	PLBPPCMMIRQ_ipd,
	PLBPPCMMRDERR_ipd,
	PLBPPCMMWRERR_ipd,
	PLBPPCMRDBTERM_ipd,
	PLBPPCMRDDACK_ipd,
	PLBPPCMRDDBUS_ipd,
	PLBPPCMRDPENDPRI_ipd,
	PLBPPCMRDPENDREQ_ipd,
	PLBPPCMRDWDADDR_ipd,
	PLBPPCMREARBITRATE_ipd,
	PLBPPCMREQPRI_ipd,
	PLBPPCMSSIZE_ipd,
	PLBPPCMTIMEOUT_ipd,
	PLBPPCMWRBTERM_ipd,
	PLBPPCMWRDACK_ipd,
	PLBPPCMWRPENDPRI_ipd,
	PLBPPCMWRPENDREQ_ipd,
	PLBPPCS0ABORT_ipd,
	PLBPPCS0ABUS_ipd,
	PLBPPCS0BE_ipd,
	PLBPPCS0BUSLOCK_ipd,
	PLBPPCS0LOCKERR_ipd,
	PLBPPCS0MASTERID_ipd,
	PLBPPCS0MSIZE_ipd,
	PLBPPCS0PAVALID_ipd,
	PLBPPCS0RDBURST_ipd,
	PLBPPCS0RDPENDPRI_ipd,
	PLBPPCS0RDPENDREQ_ipd,
	PLBPPCS0RDPRIM_ipd,
	PLBPPCS0REQPRI_ipd,
	PLBPPCS0RNW_ipd,
	PLBPPCS0SAVALID_ipd,
	PLBPPCS0SIZE_ipd,
	PLBPPCS0TATTRIBUTE_ipd,
	PLBPPCS0TYPE_ipd,
	PLBPPCS0UABUS_ipd,
	PLBPPCS0WRBURST_ipd,
	PLBPPCS0WRDBUS_ipd,
	PLBPPCS0WRPENDPRI_ipd,
	PLBPPCS0WRPENDREQ_ipd,
	PLBPPCS0WRPRIM_ipd,
	PLBPPCS1ABORT_ipd,
	PLBPPCS1ABUS_ipd,
	PLBPPCS1BE_ipd,
	PLBPPCS1BUSLOCK_ipd,
	PLBPPCS1LOCKERR_ipd,
	PLBPPCS1MASTERID_ipd,
	PLBPPCS1MSIZE_ipd,
	PLBPPCS1PAVALID_ipd,
	PLBPPCS1RDBURST_ipd,
	PLBPPCS1RDPENDPRI_ipd,
	PLBPPCS1RDPENDREQ_ipd,
	PLBPPCS1RDPRIM_ipd,
	PLBPPCS1REQPRI_ipd,
	PLBPPCS1RNW_ipd,
	PLBPPCS1SAVALID_ipd,
	PLBPPCS1SIZE_ipd,
	PLBPPCS1TATTRIBUTE_ipd,
	PLBPPCS1TYPE_ipd,
	PLBPPCS1UABUS_ipd,
	PLBPPCS1WRBURST_ipd,
	PLBPPCS1WRDBUS_ipd,
	PLBPPCS1WRPENDPRI_ipd,
	PLBPPCS1WRPENDREQ_ipd,
	PLBPPCS1WRPRIM_ipd,
	RSTC440RESETCHIP_ipd,
	RSTC440RESETCORE_ipd,
	RSTC440RESETSYSTEM_ipd,
	TIEC440DCURDLDCACHEPLBPRIO_ipd,
	TIEC440DCURDNONCACHEPLBPRIO_ipd,
	TIEC440DCURDTOUCHPLBPRIO_ipd,
	TIEC440DCURDURGENTPLBPRIO_ipd,
	TIEC440DCUWRFLUSHPLBPRIO_ipd,
	TIEC440DCUWRSTOREPLBPRIO_ipd,
	TIEC440DCUWRURGENTPLBPRIO_ipd,
	TIEC440ENDIANRESET_ipd,
	TIEC440ERPNRESET_ipd,
	TIEC440ICURDFETCHPLBPRIO_ipd,
	TIEC440ICURDSPECPLBPRIO_ipd,
	TIEC440ICURDTOUCHPLBPRIO_ipd,
	TIEC440PIR_ipd,
	TIEC440PVR_ipd,
	TIEC440USERRESET_ipd,
	TIEDCRBASEADDR_ipd,
	TRCC440TRACEDISABLE_ipd,
	TRCC440TRIGGEREVENTIN_ipd;

	end process TIMING;


end PPC440_V;
